PK
     `_[�X�,�  ,�     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_0":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_1":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_2":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_3":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_5":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6":["pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0"],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_7":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_8":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_9":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_10":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_11":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_12":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_13":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_14":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_15":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_16":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_17":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_18":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_19":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_20":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_21":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_22":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_23":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_24":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_25":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_26":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_27":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28":["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1"],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_29":["pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_1"],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_30":[],"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_31":[],"pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0":["pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0"],"pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1":["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28"],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_0":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0":["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0","pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_0"],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_1":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_1":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_2":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_2":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_3":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_3":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_4":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_4":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_5":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_5":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_6":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_6":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_7":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_7":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_8":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_8":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_9":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_9":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_10":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_10":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_11":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_11":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_12":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_12":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_13":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_13":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_14":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_14":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_15":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_15":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_16":[],"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_16":[],"pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_0":["pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0"],"pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_1":["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_29"]},"pin_to_color":{"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_0":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_1":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_2":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_3":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_5":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6":"#91D0CB","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_7":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_8":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_9":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_10":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_11":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_12":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_13":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_14":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_15":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_16":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_17":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_18":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_19":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_20":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_21":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_22":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_23":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_24":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_25":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_26":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_27":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28":"#6A826C","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_29":"#007DB5","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_30":"#000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_31":"#000000","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0":"#91D0CB","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1":"#6A826C","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_0":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0":"#91D0CB","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_1":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_1":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_2":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_2":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_3":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_3":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_4":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_4":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_5":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_5":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_6":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_6":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_7":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_7":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_8":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_8":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_9":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_9":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_10":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_10":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_11":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_11":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_12":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_12":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_13":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_13":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_14":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_14":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_15":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_15":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_16":"#000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_16":"#000000","pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_0":"#91D0CB","pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_1":"#007DB5"},"pin_to_state":{"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_0":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_1":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_2":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_3":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_5":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_7":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_8":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_9":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_10":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_11":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_12":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_13":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_14":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_15":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_16":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_17":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_18":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_19":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_20":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_21":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_22":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_23":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_24":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_25":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_26":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_27":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_29":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_30":"neutral","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_31":"neutral","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0":"neutral","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_0":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_1":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_1":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_2":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_2":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_3":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_3":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_4":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_4":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_5":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_5":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_6":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_6":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_7":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_7":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_8":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_8":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_9":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_9":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_10":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_10":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_11":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_11":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_12":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_12":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_13":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_13":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_14":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_14":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_15":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_15":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_16":"neutral","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_16":"neutral","pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_0":"neutral","pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_1":"neutral"},"next_color_idx":11,"wires_placed_in_order":[["pin-type-component_c06f5b37-fc3e-4595-b10f-4b7c1a02cd1a_0","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_7"],["pin-type-component_c06f5b37-fc3e-4595-b10f-4b7c1a02cd1a_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6"],["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6","pin-type-component_21aad173-aab7-47af-8937-bb85f96b90d7_0"],["pin-type-component_21aad173-aab7-47af-8937-bb85f96b90d7_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4"],["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4"],["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6"],["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0"],["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4"],["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_5"],["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4"],["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6"],["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0"],["pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0"],["pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_29"],["pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0","pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_0"],["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28"],["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_c06f5b37-fc3e-4595-b10f-4b7c1a02cd1a_0","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_7"]]],[[],[["pin-type-component_c06f5b37-fc3e-4595-b10f-4b7c1a02cd1a_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6"]]],[[],[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6","pin-type-component_21aad173-aab7-47af-8937-bb85f96b90d7_0"]]],[[],[["pin-type-component_21aad173-aab7-47af-8937-bb85f96b90d7_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4"]]],[[["pin-type-component_21aad173-aab7-47af-8937-bb85f96b90d7_0","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6"]],[]],[[["pin-type-component_21aad173-aab7-47af-8937-bb85f96b90d7_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4"]],[]],[[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6","pin-type-component_c06f5b37-fc3e-4595-b10f-4b7c1a02cd1a_1"]],[]],[[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_7","pin-type-component_c06f5b37-fc3e-4595-b10f-4b7c1a02cd1a_0"]],[]],[[],[["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4"]]],[[],[["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6"]]],[[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0"]],[]],[[],[["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0"]]],[[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1"]],[]],[[["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1"]],[]],[[],[["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4"]]],[[],[["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_5"]]],[[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0"]],[]],[[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_5","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1"]],[]],[[],[["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4"]]],[[],[["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6"]]],[[],[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0"]]],[[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0"]],[]],[[],[["pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0"]]],[[],[["pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_29"]]],[[],[["pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0","pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_0"]]],[[],[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28"]]],[[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4"]],[]],[[["pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1"]],[]],[[],[["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_0":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_1":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_2":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_3":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_4":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_5":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6":"0000000000000001","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_7":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_8":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_9":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_10":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_11":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_12":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_13":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_14":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_15":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_16":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_17":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_18":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_19":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_20":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_21":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_22":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_23":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_24":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_25":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_26":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_27":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28":"0000000000000000","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_29":"0000000000000002","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_30":"_","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_31":"_","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0":"0000000000000001","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1":"0000000000000000","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_0":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0":"0000000000000001","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_1":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_1":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_2":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_2":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_3":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_3":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_4":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_4":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_5":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_5":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_6":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_6":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_7":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_7":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_8":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_8":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_9":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_9":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_10":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_10":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_11":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_11":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_12":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_12":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_13":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_13":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_14":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_14":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_15":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_15":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_0_16":"_","pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_16":"_","pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_0":"0000000000000001","pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_1":"0000000000000002"},"component_id_to_pins":{"4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"8d917703-7309-40b5-92e7-4ad90a04ee5c":["0","1"],"5d364937-28f4-4ac1-9ce9-88b28ab8f411":["0","1"]},"uid_to_net":{"_":[],"0000000000000001":["pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6","pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0","pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_0"],"0000000000000002":["pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_29"],"0000000000000000":["pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1","pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28"]},"uid_to_text_label":{"0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000000":"Net 0"},"all_breadboard_info_list":["6dc8c187-74d0-473a-92ce-46ee1acaf8dd_17_2_False_505_535_up"],"breadboard_info_list":["6dc8c187-74d0-473a-92ce-46ee1acaf8dd_17_2_False_505_535_up"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[651.25,252.5],"typeId":"b269da49-8c00-4ebb-bd25-5859ea0c7cad","componentVersion":9,"instanceId":"4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44","orientation":"up","circleData":[[632.5,395],[647.5,395],[662.5,395],[677.5,395],[692.5,395],[707.5,395],[722.5,395],[737.5,395],[767.5,395],[782.5,395],[797.5,395],[812.5,395],[827.5,395],[842.5,395],[578.5,110],[593.5,110],[608.5,110],[623.5,110],[638.5,110],[653.5,110],[668.5,110],[683.5,110],[698.5,110],[713.5,110],[737.5,110],[752.5,110],[767.5,110],[782.5,110],[797.5,110],[812.5,110],[827.5,110],[842.5,110]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"3c7d2cea-7402-404e-a999-9e412705ecbc\",\"explorerHtmlId\":\"4b80aea5-44e1-4fad-a932-fe8fbd1d33b2\",\"nameHtmlId\":\"c1c471ee-6d48-42ea-837e-705af42b78aa\",\"nameInputHtmlId\":\"b279b2cc-2f2e-46a7-bae8-f6b9a233c384\",\"explorerChildHtmlId\":\"05b44ea5-1c8f-4b01-9962-f9d302a45494\",\"explorerCarrotOpenHtmlId\":\"db67ec27-7a67-4e1b-a338-2dc0ebd27123\",\"explorerCarrotClosedHtmlId\":\"d8512071-9515-46b9-ae00-97eecf4ddcd6\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},1,1100,file,{\"name\":\"sketch.ino\",\"id\":\"a0074415-63f7-4f59-920e-8ca1e1dc6f44\",\"explorerHtmlId\":\"6e8e0e1e-6c51-4861-bbf3-3d235e0462fd\",\"nameHtmlId\":\"e3d3351e-37f8-4c54-a4f1-239f80422ba4\",\"nameInputHtmlId\":\"f494cd71-e060-4966-8497-28c57457ce27\",\"code\":\"/*\\n * This Arduino sketch controls two LEDs connected to an Arduino UNO.\\n * The green LED is always on, powered directly from the 5V pin.\\n * The red LED is connected to digital pin D2 and will blink on and off\\n * every 1000 milliseconds (1 second).\\n */\\n\\nconst int redLEDPin = 2; // Pin connected to the red LED anode\\nconst int greenLEDPin = 3; // Pin connected to the red LED anode\\n\\nvoid setup() {\\n  // Initialize the red LED pin as an output\\n  pinMode(redLEDPin, OUTPUT);\\n  pinMode(greenLEDPin, OUTPUT);\\n}\\n\\nvoid loop() {\\n  // Turn the red LED on\\n  digitalWrite(redLEDPin, HIGH);\\n  digitalWrite(greenLEDPin, LOW);\\n  // Wait for 1000 milliseconds (1 second)\\n  delay(1000);\\n  // Turn the red LED off\\n  digitalWrite(redLEDPin, LOW);\\n  digitalWrite(greenLEDPin, HIGH);\\n  // Wait for 1000 milliseconds (1 second)\\n  delay(1000);\\n}\\n//\"},0,","codeLabelPosition":[651.25,95],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[882.5000245,532.5000245],"typeId":"a70bb5a8-99ed-4f1b-882e-eac0873b75ef","componentVersion":5,"instanceId":"8d917703-7309-40b5-92e7-4ad90a04ee5c","orientation":"up","circleData":[[872.5,575],[895.761385,574.8720905]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[880.0478665,622.202999],"typeId":"5f0a7f7f-5908-4e39-94d8-2714a0462581","componentVersion":2,"instanceId":"5d364937-28f4-4ac1-9ce9-88b28ab8f411","orientation":"up","circleData":[[872.5,650],[887.5,650]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"85.00000","left":"420.00000","width":"522.50005","height":"704.50000","x":"420.00000","y":"85.00000"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0\",\"endPinId\":\"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0_0\",\"rawEndPinId\":\"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"572.5000000000_545.0000000000\\\",\\\"572.5000000000_425.0000000000\\\",\\\"722.5000000000_425.0000000000\\\",\\\"722.5000000000_395.0000000000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0\",\"endPinId\":\"pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0_1\",\"rawEndPinId\":\"pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"587.5000000000_545.0000000000\\\",\\\"587.5000000000_485.0000000000\\\",\\\"872.5000000000_485.0000000000\\\",\\\"872.5000000000_575.0000000000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-breadboard_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0\",\"endPinId\":\"pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_6dc8c187-74d0-473a-92ce-46ee1acaf8dd_1_0_2\",\"rawEndPinId\":\"pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_545.0000000000\\\",\\\"602.5000000000_620.0000000000\\\",\\\"872.5000000000_620.0000000000\\\",\\\"872.5000000000_650.0000000000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_29\",\"endPinId\":\"pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_1\",\"rawStartPinId\":\"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_29\",\"rawEndPinId\":\"pin-type-component_5d364937-28f4-4ac1-9ce9-88b28ab8f411_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_110.0000000000\\\",\\\"812.5000000000_80.0000000000\\\",\\\"407.5000000000_80.0000000000\\\",\\\"407.5000000000_680.0000000000\\\",\\\"887.5000000000_680.0000000000\\\",\\\"887.5000000000_650.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28\",\"endPinId\":\"pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1\",\"rawStartPinId\":\"pin-type-component_4a14b8c6-4ff7-423d-a2f7-8e216e0a6c44_28\",\"rawEndPinId\":\"pin-type-component_8d917703-7309-40b5-92e7-4ad90a04ee5c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_110.0000000000\\\",\\\"797.5000000000_80.0000000000\\\",\\\"407.5000000000_80.0000000000\\\",\\\"407.5000000000_605.0000000000\\\",\\\"895.7613850000_605.0000000000\\\",\\\"895.7613850000_574.8720905000\\\"]}\"}"],"projectDescription":""}PK
     `_[               jsons/PK
     `_[1G��  �     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino UNO","category":["User Defined"],"userDefined":true,"id":"b269da49-8c00-4ebb-bd25-5859ea0c7cad","subtypeDescription":"","subtypePic":"e30496d1-6e1c-40fa-a66f-2add70ecdc94.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"a7fde0f7-2836-4f0c-aad0-66dcccec46ff.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":9,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"LED Two Pin (Green)","category":["User Defined"],"id":"a70bb5a8-99ed-4f1b-882e-eac0873b75ef","componentVersion":5,"userDefined":true,"subtypeDescription":"","subtypePic":"f9728bc6-2422-4ead-9082-90351081a874.png","iconPic":"9ba3df0f-d630-43f7-8169-617793654d93.png","hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/3749fe76-cef7-4b42-9f27-525b8a44301e.svg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"8.33333","pins":[{"uniquePinIdString":"0","positionMil":"266.66667,133.33333","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"421.74257,134.18606","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"LED Two Pin (Red)","category":["User Defined"],"id":"5f0a7f7f-5908-4e39-94d8-2714a0462581","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"3d0a314b-f708-4b2c-819f-35c414b123ec.png","iconPic":"6608fa58-7afa-4488-b64c-2b761d69d6bd.png","hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/a9e23d57-c0ac-465e-ae7a-a15cecbcb7b3.svg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"4.24452","numDisplayRows":"5.30565","pins":[{"uniquePinIdString":"0","positionMil":"161.90689,79.96916","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"261.90689,79.96916","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[],"propertiesV2":[]}]}PK
     `_[               images/PK
     `_[�R�W�  W�  /   images/e30496d1-6e1c-40fa-a66f-2add70ecdc94.png�PNG

   IHDR  u  v   ��:   	pHYs  �  ��+  �	IDATx��	�ם�����w�}!��l��Zhz��@?aK3�`l���-Ü1���vws�c�w������=��-,��lt��#��%K��� �ElE-Ԟ9�ݪ�����̈��ܾ�9A%��q#n�ȼ_��"!�fs]uD��$�\B�0$R+�B!��� &�t���4H�BQ�&�뿿6�m��#�B!$71��_�yd�䪰��s˚�u5��NC��-�B!���&��E��]S($7	!�B!$/�UaGQ� �7玕�%�7��t����˒i�(���F��C��B!�B��EaGQ��u[7a�����������!y�ђiF�����!�B!�&ׄE��l��emM��8If��?�J���2)K��̙3�ih�kB!�B�p䒰��s@u$��X^e�������r!�B!�&W�E�A� yD!�B!Ğ\vu`�KB!�B
�lvu)R���B!�B)H�Y�Q�R �b�4I(z4����±ȼP(6Mb���hB!���d������gL�ۧ���ή��^7n�DB}���'�;"��|���)*�Hqq��_����}�Cr%�$���';e��a6m�/J�l�V�,7D�Z�Kk�B!��Ad����������'��s/^��󘢢"Yq�d���������_:}2�D�\_(����uMN?۵u��.�-��-��77�B�w�B!��6aGQGH����6�>�-^���u��f�Κ"%�ֈ�,����3�z�����v�.��]�X���vٮ���@6	;�:B�XL��D�~w�>Ow�u]s��ڪG67�%�h|y9��1���2���ns����,��v�.�e�fڪG�G��)�R�zA��pϰ��S��]��o���ϧ��lvu��8t-}х�İqsi���u;+ݼ�(nr#�!�B�lvu��0qA��?A���B!d(�vu��(���˥�:+vU�ln�H�gB!�B�@�2�6E!9JT|��K�b�<�uk:�S����̮(U���]��v�n�+�Ѩ���z��P($�)��a�l���n.@QG�����S���������:P^^������%_n�leڞX�3S��F7��ܺa����tww�},��%2r���8d�l��]/���������%W�^M{_�pXƎ���e�l���n.@QG���z�����ܬD��Ç���9������v�T��0A*jj���Zjkk��#���m��l]�[�ym(~����EZZ�?&ҙ�ab6v�X�%����]��v����D"ERQQ�քTODQw5��(�e�l7�vs�� ����Ւ
��w�Tg��@̝?^.�=+'�~[�����bn�!�ʌ�!��%1��?�=��5^�?�W�1y�x]>n�T]3C��~���4IF��D^&�(��yw����\����Q$<�ǁ:v5�lݒNҔt&hzb�/xL��.�e�l��v�"�	�y"�v�.���l&�Άx�\B̝<|X>nj��C��Q#��j���s����i@��a)���R,��v� o��5)�6M�/�s�6w��3&���Hn�h(�(�C��Y����<1c�l��ݠ��
7R/&�l����t �Έ�n��s{�Jǁ�2�s��e�q�t:��]�q�`�.�H穓����rd�T��?�/2�����^�3���J$K�G���D��>Jy�Oz�'3��v�.����^�p!���k��Γ�(�e�l7?�O~�qŕ+W佷ޒ#��i55Rk��+��K�"�G�ʸ��"i;}J�ܺE.�志ًɄ	�8 &M�E �f�#[�xQ���=�'m^�M�]��v�n����J����a�l���uDA���.W^��\?�^�;&}==��qWq�ʱ�~"��2e�!�a�I/a�͐�#�B!$#P�%�~�{�D��'�*�����(~ �$Y_V&�엽O=%���i�K�h8�$Y�f���B!$cP�8����C`���ʩS��[Ɉ�"�|��4��?ɟ��*��B!����Y.�񆴿�[�PV*�t-�.��7������+�ň$��7��/a=K��B!�d��Y.O��_�5u�r���(nP®�Hξ���;�]'�.^���B!�BR���@���;;��Z���C�
���YR"o�h�L�9S&N�*Ğ�"��.ٕ3/�pB!���AQW����_K�'�'��Ύ����G�R��.����e��մ�B!��"uHgg�m�\S[#�?�P��;�,���W_�O�/�q�&	���e��θt�B!�d������Rc���u��Rˈ����K�2��P!Y(�B!$cP��?u�|~�ti��J���Q5���"= hj��UUr��i�&`�+�D�Hӯ������L��,P�n��J��3fL���W�]��v�n����K�������]��E�fu2��J���P���}\\/;O������ ӥ�v���r���y�g��4!�ڪG6/o�޺��E�^�g���r�5�8�L{{�tu%@�v�.�e�^���\.X���gp�8��v�nf��F(�
���pD:._�l�(Vֺ�R�% SB*+D�AC�;�Ĭ�������6�4��v�.��8��c�:�\ii���vB�v�.�M��l�����x��T��I˙3���6�غO��!��BrO��Ӻ��;���^����t��vb����g\�.�e�l�i�^�v"�q;!e�l���n6CQW`t��H��2^�`8"�R�t�!�)���$��uk6ׅB�-n?�DdĈiM�4�b��b)�5�]��vٮ�v�"�,�iND5zB��ő�]��~�� E]��z�Ttg���7l�E�p]tw&c�j��ӱ�Iww�\�xѓ����]��v�h�+P����]��v�����("��^�v`�#��pcţ�^��}A�1i\�5��#���Yа]��v�n������]��v�:BrXʊ��f�Bٺ�9�6Q� 5�$�B!YE]�Q\��<LK]J�BrSM$������+����M�B!�B�%7f����ha�����\1�r	!�BH�AQW`�"ER\^.�L�:MuN����z��7�>�5�Y)��fs�@R�1tg&�T�p,�u�|��X�j��t`�l��]?h�%o���n��׋�]����+0FL�,��[q�X_�d#�XLjg��X�B����[����ۿ��)���:t!%覊ϼxe�d��v�.��/�z�]����f#uF̈́	r�w���L����b�!���O��;(��q�JL���}�3�x;5/�D��pmb�B!��E]�1a�l��g�IyMMV�:�>c�<w���I���"y*��&	E�FCrԼ]8�g��i��p����B!$7�����m���Ei�L^�{��U��kJ++���LF������6 �:�1�~�mB�C	<cQ�톼9 �Ƙ2Kgϐ9F�׻���!�BH�������jI���U����<o�Mz����/۬u=��9g���ds&���|Ff:���[�çdE�.�ґ��M����>-�&��i#���xE���D_?(�9x>�BH!BQW�\w���jӯ�v�Ȭutݱ�|�s�B����R���2�<�z�{fLTbo�S�$W�3�g�ßW�BN8��M���E�e��?S�B!�E]+��[�T"}�Uֺ�hTb�2��[��lc��k	���n����D�]r�52��F�_j�\ �®�!;��h�{v�.P�,��}�8�K�I�/��Vgg�kt�⵪���l�

����%K�x]F�-��@�A��Jw���BH62e�k�@�-���z�{��qawǌ��#D,q�"��Ϥ�CއuNY�6|Y�ϽV���wBH*`+���&�1���
� ���P�6[�*ʔ�0�	��xcz�O^�J˳>�-/�����KnW}��e�p�X�q�k������~5h}���Xi��l|�ׁ=PjZ�����X~�l|��� ���E���1�����u_f�3����(�
X����"���[R9r��_t^��+����z捴����,%]W��Gwi�|0sQ��6��(ǧޜ��%�W��^�p4�z�N�M���G�NT�~�0yHֶ��m��#)�]z��������k�'��k=Ld1�����'�j�j�O���H��bw�R��8�lu)Ʊ�_^?ŗɽ�O ��O��BM|�=����^-00&������t�w='ZLڡ�����n1���O��y|��ϸ/���>�p6�86W&~��@���-R�~��v����𙄢����t�����d����~Uz:;?�]�4]W8"��o�F��:���v�o�-�zE��ًmw䅣�o*�n���������u���B�_k�>��>�)�ښɤг��W���	��ǰ�a��ɒ�Ƹ�$�1�!��ˣ���6_�E�_YA,�Řઉ��>�q�jf���)�t��z��p]О��Ax��%���7=̖;e�B�|?yٓv��8�����x�u�/�PlZ��|�=��z|zu��f��M7��3����7c	�m���~�}�o,)�
�������o�������Gv}}�J�����/}�+a���Rv^�����RЙ���Ϟ��o��ՙ�x��#i��%z�ݐ�A���uB[i�� �u�fr�uz��, �yjV'c�z�����gF	��L�1m0�_Y��0��x鎨,9F��1��A�d��m��7�S��w�����ǈ�hA����B���ĸW���Ό���z}���8?�+������1lN��7�74������񷖢������kk�7��]�0i�\9y*0a��^����ZXi�	;��N��!�4��������M�T� ����g_2<tC
�̮ts���~���νmZ}� k!���D�ڮ~�~0�����X�(7[���t�u7��>��
��ۆ��n�����z��A�,fk�c|`���S�l�����_��,�;�/�+�)T���3��H���.�ʊ�"��%6���#2j�t�w_T	���������ꀅ�S_]-��Y|I���&���];a秠ӄ� +�<*s�ޗ�����Dx�Y�nH���VgGܽ�C�:e�o��,c⌶!�!Lp]1��>�߫k�����/�ԡ-sL�H��7Zܩ{��)����DL�7������G�[Q�^N�16�����\@�v1Np~]/|��G�Xt�N�PI_�v���9�c:p�xy��ݍƘ�k��J������Qň��kE?$Ľ�,ۖ�E}}���7(��n�?l����q;e�\�xї�)���t�E�/���~#-t>ⷰ�X�]P횅]�����?��>$O	
L�Ryr�I�����ܐ *%f��ۧvGN���ަ�_b���ya�:L�0q�rB�bhD�.�ؿ)_Z2H8@X��DN]+�
�Mu �cU�K��Ճ��X�u��	�����"���@�^�D?\~=��y@ kwD�}���xy�hGd�wf/���OQ�Ǹ�A�-��a��Ȭ�V{�Pԑ8�c�Ȣ��[�����+R?m���?�I���tG���Iф�x�7T{��m2a�A[�~]�� ۅ��-*����t�vOO�1��(k�%p�n���S�$;h
�IM�&A��K�i�x=�18`��dj�O.Ov�Ƥ�j��Ѽy_&&���t	
s������o.��N��^�� ��NFa��^6m���!~��g��D��8�y����>��I��'�;�vPI��3u�Eb��X�ZN<(��~Jjjk�j�h��N��h,&��R���J����	�t��!�ۓ�v+�.*���%�,(7@��p���+AYhnHzb��?0Q�F�vu�3��`"�[��,�WɅI�~=Â3���A��*�@z�D����&���_�gɚl���������	���w��_���Dj��$�"ᆸ�2�X��D.��=��9����ɍ���#�D&k��5%Yjo�5�y:���2i��㔂�쎘�:k׻�y�,�B
�� �{��}�8i�Ln�YW+������w�?.��|"��쑳o�!��=RZ^.��s��q=Ʊ����װʕ�+�fϑk?�X��e�HD�r�t�K��8���}pD޾|�>���rdu1�KL�G�:����x=�/D7$�~aԓc�V��l��˥�BH栨�������'��/")ӢN���y��+r��u��Yi�l�7WTT$+n�,��1VUU%����y+��g���d�	��KW���.9�Ijc6�v��,���fx�r��nHΞk��v��Ep�q>p9��h��=�p�U�.�[
��5�t�h?\�
�)��_I6�1g�h��ٕV�F,����������,�q2����:�f��m�GTIEE�||�^�@е�uH4���Z�(�ힱo�V��mF��Ew.��+���Kn�O;�a-,R�<~�]�`�D9x��,���\�e0��ص�����$;�|��6m�<����E!��1#�K������ܦ���H�(l�;8وj�V��n������2�&d*�?��]3�^|CV�5O��x�lX|�<���B����`\��w�,���������8Yy�Lyp�̂'��oճ/I!pǌI�/Ɠ�u]�`b��{���d��7��|����g��9���A�B���ۭ�����B��v�]� qn�Ə���L��g��>,���55�"�&����Sn��+WL=N �
a���)#j��X¢Y������T�>&�:B!y���a�T�L��g�������d�xϝ_�B'�t��fA�?����X�w<�$���[��:B)0�����<����i͸��g��up3��E�aJ}���z��#��{���8)�����վ��½u��I�u���JQG!�NL���7('T�s;2����	q��!$�8p���\aÀU%(��q�J���B�/`��=a��{_�s��:x�s7Ld����e�=w%�,`��G(�)p.\h�ʲ�5��L-m���nSK̻vۤ�|p��)˥��5/�5똝�J�������������l7V��o�ض�m!�b� �N\nl�[h�P����Ҋ_n��]6{��8[���<NNCQGH��'����G"��_���M���;���.�]p>9�*�	^���t�ty�ݏ���L�k��-�J���khX���E'�@E���g�(�qR(�k�vi�O7�U?~I��_1��.��HP�ȏ��H~}�tt'/��S�ejU�oA��G_> �p�X�I�?u�W�[%�X,�p�k�����O����n_��n$q�ӧ���{떑�v�G�{��A`��(~nqY(q@�SP`]̚�GOv�"�]��B'�~���.���e�/���3��.5ur�r�ZR�����b!��F�3�BD���	����3����v���ue��'!��������/b�T�������?�ӌ��N��iWM�{l{u��B1���R��Iv�/\+\�c�z����B'H�s���Źٹ?��+�cϿ��1������E!�d *X�t����)�����+��%���.7�p�l�_s{:���맨���8b`�we�1a����@d {��	������+�qR(�q�K7$�5?)!g���B2�v}��!������z�WE��K��@�!^.YLl�v�|!���ڤ*��Z�nj�6N
�|���u�P�BH�����
��Ec�K&�����VAa�6��a�öX�0%=��b�L������m��84\�$�������)))�p
	C���3�t�d-���\O������:gwV�"R�9
���2�&��{�-�T*�L�}����M!$(겔�HD"���]6��P(�����z締C��;��a&���pE����e�C�Tbě�dm���fApB�'(겔ʲR)-��������d�7i�<�ٛ��B��%����H��!vo�O^��Y/����!�;��:��U&8��"��(겔_:#��?����.I6p��]	LB�� ~A�,�5����q1�R*���z�3o:p����!�!҈�JG!�E]����u��6N�td�Ő� �5K�u�u��%IQ ���	qg�m������r�j�Q��R��[f����p�BH!AQG!��#v�jAǯ�
��t�<:���Æ�d%(�|۷��MQG!y	E!�d��[�Mi;���f����B����T̘('.�����(��<}�qu�������8S�BH�$%��^OV�ض��
<��{��];0��Dۄ����	�
�W{��vU=X�4_C(��L���	�GL�d̮U��X̟A�nX��y�`���i?����X�q;G���m�,38�T���"�F݀�����	�VӇǅ�6��!I������ yPV3h/ȶ	!�I&��CVg�}b|�Y��`���w6�uy���0n(��^�}�qȓ�i�dJOO�yd���¯�L>q5�}@�$V7�T�h�D���"� x �3N�}Z��$Fy��W��{�V���>��3�Y��2�6!��Ȕ�B���0�x�6����7�E]� +/n2u��ȸ����y��3�Aԩ�}	�^B��%e�3X��%�����G��.�����j)��	!�E&�~Ga�H�/��bN���|����Ж8�Y��MR� _��B��{?f�a��o�b���e�B�V2%�0�ł��{(��S	����)E]�I�6��z�UΘt��͈xB�3�?>�u#�OB�q2)�0'���]�Q�Z��U���k���u�ʠw��x�+�a��l>�M��u��;'n<q���..O%o�I��m��t�
���po�>�}ń(�Br�L�+�0�p�[���y!��E]��ڌ��p9�D)�9�?�3��e����n�n"�=k�b&| ���a�����U�"D�'��KdR\��Ƃ��AY7����i<ɘ�曰���C��/1�a)�ൖH5�h�Qt�X���g��F'3�%�c��
��`���	!��
��+/1']Q�7m~71n���@5�uyN<5�W���v��TQ����e7�Nɞ�O?����,��?�_n���Cr�\3���`�Vp�<�wu�Br�D�J�՜��q��06����:Y>z�P�9�Ϊ��-���������TC��cIC��N�n�tC�NS�����RQ�����}���M��*��p�'��BH��J��-fڃ�A���aP�--� ����R��ytd�?I�!VzEƗ�%�� ƍ�B��%��q�<��a�k'֍�U�@�;�S#���?qi��K����B!$U2i1üT%�3�=j�nr��3D�.��C���������@Ow׵�����	M��e�� �7���x��͙(�%�����,���칋�օBl�B!�ȴ�L�+ю����_�f>CQ��p����8�$&l��R�
J�J�.a鸎��!�BH�i��99�O3�:B!�BI�LY�̞d�J�e����:B!�B��m1�xӮ�?|!���c�^�����ˢ��E!΅mRY>8�㔉����*�W;�.!�B��L��`�����.�X �X���7|r�U:;:$bI���t�ty�ݏ�Ӈ���.!�R(d�b�6��vj�Os��|�������V���J,I�͵ӧ��ߟd����P`2kEե|��!$����5y��bҌڱe	1>o�Bm�<,$�&��,�zbng���I�Sk���c���=o�6����Xp�Ȥh�}>�����.�4o���z���.C7��m�r��s��H&�Le�b��2������#u�(��|f�ZZ��b�*�0߸�v%2�Ց�b�f=i��b!`Y+��Q��DYqL9J$�ʛ�O7�%��˄�2&���p ��b� �͢"m`тQogm��^��˷I��K�%��1�'�wӇ�n����7�������|���%��#�B� z��Č1	Od1�d��:�HC.��v"
� �����Tn��T�G_����a����)���1���1�zhf�����?���
s&����Uj�J���y���e���&+n�)e�E�7����E�3�q*V\��������	�ځ���{+_k�Q�B!�dL��.�=n!�COJMԭ�hݢ�_eU���@(b_N\��W����O��2-�v�?�D��?&�X�Qh�� u�z[��,� ��D.�A1��Fv��Wj�J���Dyp�Ly��)ٶg��>xX�_9��0�^�tve�Z�)T<�3�J�~���4u��!ݥR~5�:,}E�i���^J��$��x���%v1fLL!d�D[��(ڃ0H���#�c׮�f7MXӴ�(�����f�mq܉b����	�K��`a,Y���Q����P,rpfLTKKg���"�'���[����a�S>�c����}���93u��!�\$��h���@��*��#3nS��l��irz�ra�t���I8�h���5��w!��;���范N�qfں�8>�
��]
{��X̠��&�ɹ��iˡ�J*17`�3[⬨�+Kn�[q��LZ��P;06��٧��x�}��1c���k�,1D�t+��%��|���� �"(1��.�]�:@QGH����Ł,:�t�Vǧެ^w�T��7�O�;s���%����٦��ٲ�J��d(��I��]0X�Rbb�Nh���c��N��ר~���cj���""�1b=D���t��\���:+����Ձ?��)�� �~��[ԙ�w�E!y���*�j�NX!�(�!~2�,��d�.�~�}C�4`1�;��D�, � �pf7Ns{U�`��=s�%�S�K$ˀ���x�G(��s�X����'��vt�?��PI>�qS5�P� MW��AŨmzz��x]:����tK�uG���巆�7�s��S���[�^o�$S�dsL�S ��A�	�f��k�N�J�'���o fk������X�%�WZVv�'��.\M�~e\HH0��rLN�� �V2A�W��+?�!�OT"c�9\9��0�5i��-�4��3����D�Xt&�t�� .�IڡV�׃�Cܟ!�e�4.�Y1���w0����O��P(T�F�4S���y���|�d9�`%��z]"�O+h#��p��7&���,%]W��2\"K��6���������^I[�9i�BR�L� K�X*�	� FH%4�ǯ�׫Zl)�K��&J��\faf=�qX��ݢ3]ډ�e邔�� Z��x"p�2Q|B*B�Jz�*��N�X��awp�_!�d���}��)oߐ��I��$n�ü���}�#!���y��Úf�P�tnu�$�W��֤,��;W����ʄE���U���#�B!���$�ʹ!Obֲ��$w��#�B!���S�}@��J�W&PV:S�ARP�B!��@�k��X]eIa@QG!�B!9E!�8S�kdʈ!�B
���˕<+|NQG!̜	�e��{���D!��B����t�sy%�&N�x5g� *++�kkk�������B�Pv<����BHA1{�(y���dճ/I�@K!y��o=�
�Z��Qd��^Z��>���Mdl���Z�A�2c���`��/�ׇC6�-/�5h�(���梴���~����ˊ�v�RG!������_�|����D/�2s��	�a�u��z��^�����,kafʹ�m��P��r�O^V�v>�y����a�;��\�k��/��lqw<��1u�B
��Br��-�-R��,� DX]E�_���[��.��D�U�A��3 �O%}2>A��! ��@`BB�xj0�ԢB!��&u�`py�����Ġ��9�BDc��uS��s��B!dx(�)0�K�x�2���->�YӇ�Ӳ�Ab��2g`L!�BHr(�)0`�j����3?|A�l�D)���0�IR�hft��Y4ڶw�l%�Rq�$�B)t(�!I��S�S�E�o�Pg�T�Ol����*�bF��g�C�X��~�B!��:B
X�҉UӂLe¼�:ٸ��x"s��d���@�S%`I��G!�R�P�R`��HY��F�(��jZ}�e��.90h_�|��S�_?eP�:��B�]:�!�B)4(�)0��R�N.�o+�t;����z;�N|�*n@�ڃ��N8B!��ᡨ#��� C]8U����+�,n��A�i�I��-v(m��%�A ��9�PG)4��ר��S���s�$�r���B�N_����`��3g�hc�^O�33�c}����#B��#� �{�W�����!�l����ֺ��z8��O	D�Y*!!վL�a>N����<�d��k�h�3q�Ԕ�������!^�>)�Q�/_�p�}t��LQ��3dh?�tv��9tR	�|�#'<~�]��;��x��WdǛ��n�^6��g��;{ze���&?}�C5>w<�L�9��cϿ��ͺ~E�.��a�-3e���������^���������}j=xl������o�_o>�m��-���F�c�1c���gʉ˭������w4,S�֯xj�:v<8�~�g��Ot����r����\x���#��?,�[�z�\	�Br��U|o�z��l����<g��=i�Ng�L�T�[���v@,&+o@��S�Je������N�Pq��G$
��FGw�t��Ji�a	�'C}�=r{�a�W0y\}�<C��H*✀I*L�1��}�<cLn!dr�eF-��O���ƾ��0�Gm3DF>Z�0� v�k�!| � �c�!n��t���H��:-r ���t�s�{����o2����Ȃ�t�Ѷy=��zX�1V���m�1b�pXf��m+�c����C��1O��Ա����|�����_���*��G�|y���~*�qS��'�U�Ͼ�\m�q\xb|��1��u�B$��%]���nҵ3��"��$e*�$�ʙ��Jg�Y˛!�7�V���]��"���y�1!���K�k�&�Xc۞�s��R�������P�-ܬ�Z��*�cb�R�Q.�X �*֐��N�=�}�;�v�Nm{��59����q�և���hA��7���v�6g��ScWO��2�;�B�_�	(�!����vJ����HQ��yդ�k�L�6|�6�EJ"���o�~��l߳O�� Ŝ�'�R}ѝ+،vc���a�^�"j�,f�����x `;/�{DY~a	6�_�,^*\�l�X��} C�����"iuK��cv���p�4o�s�;���h4$�.�wʫ��&;|�YY���ߕu~@�O�;)!~BQG!9�.9�.`2z�;����j���>c镪�	R\Z+d(�
�Z�e.0	�t�]j�Mna��f� ��{,G\�0δ��������"��e�qiE�~�&�W�yQ}�f�8�M�|#�^�m����/�c��Y�#�N?X���B뵘�k� sL��c��b�������a�1AP�عUϾ�����S��Y��[�����/�ԭ|z��{�<���xL�'�W��?|AV�2k��D�b����;��*L��:B!�Ģ}���+�XL�Q'a�3�>4&5Q5�)�-䏮o^ły�v���L%w���+Y����d�!H��}���97O3D`œ��k��XQ	D��Ԑ�Xv�!T��J��uvV+�cL�^%bf������sJ�����������X�;(���ڕ�����(��P�B����Dj믑�1I)..��2���弜9sH����ȱ3%�H��bN"��@t��CJ�m��eɜ$#[��|���D��L�������E�hK�C��	I|'X�,�#�x��x���P�B��~�)�9d}U�h��>�_Ξ��L��))*�P�uwwK��I�9�_. �	��#j�4?����g�u.��̩�3�ϚIr�qL86�����H2,����鑋W����_ƷQ.��Zs6S-�N(�!��b�r��a9{r���t�!�
'�
�u��\Ǯj�m�7wL��7gd�50)��ʤ˪]vH$��u˴�$�����Y��FKQG����B�kƎ�A���������qR?+�.�4���s��</̍d(H����eu��{}�v@p_��ms���O�Bc��3Q�OBܒ����B|e��OI��c�u��T�^���1�tV�)�/�N��d_�㪷���X�襰��'�l�S�Hh�,��9C�j"��hn��Jة���e�p�5'@��Qܛ�p�EB}_�h���Ol��qW�,�$?��#����f��핎N���>ii�Pƌ����1a}�R�@D�>xDձzͦ`s"��i�;F�8��W�Ώ,�8�g�	1����b��uA����.z�
c|�S�c��2�Ȕo�@Hn7^Ǌ{Vr회k��AĹ�����B�k*++����~�\��WN{�vb+�}��E%׀0���aiy����3���c��u� ұ�+�0I�5ˋ�(~�ъ[f�b����*&�~Ʋ�Ya}�M�˼�d�b�E!��G�d┹r��>5�[J�륻�\Tu�@�/�\� `�I�M/�w��
��ҵ�Tf�ŷ�v=LG�y����>B6B,�|��܊;��ç|Y{m,�t��C��BP�m�b����k�6�	�/�K��c�I�:B!CGJ��l��!RT*�'�$��~(}�HQ$&�e��s��~�#��v���?��{�᳷)WQ7�v�l
b�
�b��7�d�n�������(����Y-�ee�neUی>I�X�5�`Q�*N�\c`��X,���p�������z��1�����B�@�8�!�p�9�N c��㇫0��z�m5&u�AB������B|�f�Jع��Q� �����6)��H(��r��8r+X0�D�[B7`��:f�n,Rv.�$I7)
&�8���M�2���Բ���dܫ�:�K�!�&�ւ֩ �c�^&��k�����9"�za�����0���N��� �-�)<�I5�	�@���k�W�߃v3HaCQG!y�ƥ�b��-�ʾ����/�����q��?�S]����hTB�L�+U��	�`����Y3�������25at
\)!x��X��8_XU~�A�B�ќo?�,�fW*���8K/ĉ���|N��s�}2k2=zU~V6X[q�ZHa4q�1�u���P�B�3�"t����¡6);s����$*�Cm��CG�����=+�b�ܸ]B��J�X��m��l��3��):#��K��v"75�o?h*M�)�Gp5u#��7^�:klU�V�L�sŽ��ӽ.���_��K�-�ΪJ
�:B�a���wjI��WE��UX�u����".O��e�-`1D���2�� ��jw�:Lt1��&ᢅ���+��"
�6���ǞE	o����+�a�M4�f�W;p�c4[1FP3.�v�n�R�g�x�JG�BQG!�XX���=&�?��L�:Q�a��붵�I&&�n,��(�48&XQ��I,چŷ�up��c`"����'R+��U�l�
. ���ڼ��eELtTɍK��Lpq@��q�
��Vu�l���y��B$}(�!�Ȏ�<��d]*@�!q�SWL=A����|tXG���qn��̻��Ä}ת/������l�3�*"�m{����J��v"�q�C���h�����b_XplڵY[�i��-j����5A�KQG!����q"\tz�\ ����%D��	���mpզW�Κ��چ1Z��\6�G�eV�Ź�춧
�ϟ��	k� �~�H��(�#��۩�����E�N����\;�.�*��z�i�CH�ˆ����E!�bb�C��N�e�t��ǉAܠ&�Y膋qD<�W�7T��o<���Ȅ	�O�V�+��o��6P�M�uy�dXE���ƣ{�i-�0n��ֺT��%La��$��B ���
[���uK	;��cN�ݖ����	�7ե��q$
v���r�� ����|g��S�~1t/�C$c�ML)������t�/�18�����S���⌱`���
�_�?-�(�!����t�b2�	0q��C;���,��aӋ�;u��:u ��*9
�]@w�3q��"��Y�L����1��W�b y�5q
\kO�Bk8w�h%��ͮJ2K���B�N�����l�v�
�򇉦������L�� ��V���N@,jk�)�x)]x�����uA~׮õ��F쵅.���+o����C�`[;�M����ݴ��,A	;�:B!d '�s$x�u�f���|����!LSu�QL���f�<%f
0
*�]�ᒉ>�+ӣ����A��ZE�3��RM��qg�bF�~���r� �E!�2�5{�p<��{�@�͙8ʳ�)�~�R����с	�q���d�Į�5�NHc��!��_������!�c����DU�.��|-5p�gG�w�vu�B��#Q�'�n�Ŝ��&�n-^&N���k�O�פrmR��9q^�Z�`�Lep�4�\�1�"��~�� �����������gm/�񡱳���"�㧰��#�BD	���M�[;ae�n�q7��gJT�9t�?���7{�?��87Ba�1�NU��i���%y�\-�r	��9�l�����3�{�Ə�uv ��J�r���cOu| �p��CY�<�K�Q�B!b��.�t~���L�MPHۭ%�0�K?�����H�X��:�Ŏ�������~Ԯ���~Ƨ��^�J]qxk��7�J�o�!�(�!�q6�Ǥ<�0ۻ~����z&�Dpp�1O�~欏Ȋ�WY���c��d�:?���͙�,f��9D.�,���uy����BqȕN�ie
�ab���@1���M'�Gkm2;V��n�]��k@������e�;l2_��hg��SH�_�L"C2����B!q`ep.�r��8����D�l����If^�[x%�(�!���ضBE��IA�)� ]��$��ɚ�U�:���	Ɔy���u1Ib�vu�BQ�:�^��{[����&b�PDz����"��lz�Kf�Ry�vhgIv���)��m:aE�.u�Ȓ��R��B"]aGQG!�8�67��0�|ͧzS�=(��a�m�>���Hn��5a���;h��5L�e4t�7���iRM�����1XDQ���KX�En��V}!����u~�U��=�N��]��\�6�#�(�!�q6�a̙��l��W���t�yX�|�)�e��L��}��a?k���).��p�3g�D�Gs.	�Ar<�CM����F�)�C8I���~�����*q@aW�vu�B�8���7wC�]�~���&��|o��M,�k�Ǆ�N5�섃X��j燨���c�G?���,jҭ]�(%D����ڸ_:)�ˤ9[&��p٥�/�;�:B!D��.t�~T> +�V)LFw<웋i�,�}��ʱā���u07k��	���_�m��֮�&�;|uw�<`�X����B qY��Qa�����s�
X��
���iҘ�)Ydq�%s�=w��Ch��hY���<�bj�X�b�L$�Y9� !�N�:��U��J�u�<�+?�����n�[�p/�f�˂ĉ���#�B������ŕ��k^΋:�+D��`R��=w���$���[f9�>մ�p���K �:^�Y½���&�i"��?�]�_ԁU�ڻ~E\ܤS�n��#��% ���K��6�O_p�\B�`D�"�x@}N��T�E!�2���f<��UWCX�y��/sU�BD����p:i�eԜ0���MYo��y���jy
�R��1�̶W���A׮s
��Y�q���@������3o���>�᳷Ƴ�"��	RH*��B@���?��a5X����k`b�{ս��`���G�DpA3'����%��;��	IV[#�J����������@H�p�m|ة��� ��&i��u�_WV�4��W�0k������v�C������6A�/�	;�:B!d <��S/�&��8�)� ��N�3pG��	��aB��J�ɂ"�oV�򖙆�IO�-�$�A�
E��Z�g����C����)p{5Ǫ�t3kj ��\��Z���f�$��]D
��E!�bt')��!W��zr���eF	�����mϥ�?��W��q"x���T��5՜��+^����[f�6Cȸ�7��;r&�,��j��s#v ���z_���n���
ƼS���E��<�$K�#����#�BL`��$f.%A�x7�.19�0��]�F��W��o �pP�@$8.�Hq?g�(%4�\���M���&c�f����\��u�E׮�L�v1vS�/k��X���ͩ�����5x�/_w�����{�1�>���N�Q�B!6����Y�@b��քl���L4a-YѸKe#t:��a��4q��x)3xx������F�i`��Z��o�FݷT���!�.Z���2��}��k���ƳٝSa��(!�L`�:7]�~��9)��XK�����j�xVaGQG!�X��w����L�1�#&�n3]��'�zB��21�,� |`�r
�t�d&��6' �k��i<�EV?�~q��e\K�?@��K����V��S1�kdWcd��h�@F�T3�&(0�����!!��XUl�����E�!DX�{ ���T��2gC�;���4��I�Y�Q�B!68����lv8�:X}��Lpa�q�7@;X\�ʊ�.�Ļ�
a�=M�lm��6�M`�k��*� B �ƣ�\!�!�>��p�*U��N4��w�\<qcm��ƥy)�����O�-�(�!�0�[9���lv�Y��v-��>��2���u�M�r%�V��Lgu+耛x)+�������	��$���c1��)�VAg�L�v�4[�܂qk%b���m]9��_nBR��BI D�]�M20��s�$e�ʄ�!�J:Y.SqC���q����D1e�g���K�A����:��"=?���7�U�}�����֮�p�����;�[�Z����:k0n����;�҉�n�:�k��̠�>��D�mY��Ld%�E!�� X'0�vc���l��Qj�dZr����(W���\� � F�Z��Fw��TeلE�1���4����������P��3�6�86�,�Nȸ9w�h[�O�1Ch�Z�eb�ly���K�Wh����$�,������J�*17`!�cJ��e�U��u�B�0@�����*�]1��ㄏ.U8���F%rp�.]�$A&�v�[���"�S�T�)��#X_��t[���y���Eg���jz����.���ע7�[�y����bH�[(�!��$�M���-3�q�'�^&	���uN�YтΩ`.1� ���ۦ���[&���nAp�x��3�?-f��t��BQG!�$!�T�f���dq��#���aW"e��*C^:V'�[A��J؁�b�w�V�]F?�}Щ��d�ѭ�e���B3p�����s�}\��7�N	]X�P� �l�@I܁q�4�3kL`�.�$?��#�"+���ݓ�(V.�TIsU�Ģ�!�V�*�J*�5
IkW�L��:p�C���H����O��(�.9�}�hA>Lܛ�I�Y\�b�"*]k��t�F�tNX�(�`�귞\�G 1b�C!E�bW��[`�k��g�^�@&��^ƒ��0Ǻ➻���\�t�A���t��#��F��[J�.I��Q7Nr������*��#fI���ɒF�TɌ�1R_\麝�!�||����Q�Q'9���Όj3$p����px%�4iX��
��(�84k/�=����5'/�w����fe���W�|��G����K�b���"�p����핮�^)�8�~%���_><u�߀����E)-�����M#MkHi�}'?��[���^^7Y6�~M��j�B�<쳮�Lm��;X��[��m�"Cȉ�$j���Z�(M?���e�vA㶦V*`�H��@y6��L�<���k��C  >�g�z/+K���V�v�V첏zJۇ��V��O�ȑ��F=k�:��Y�l?ky'$�B,&�KS,�i6��ɴP(<��	]
�M~E!��?|A��m�l\�@	���Nz��KKd��ý�'/�t�Ģ�r���?wD��kd�\�������-쐒<l0��uֆb���9�G?0�'�.qh_gI�˞�����x�r��N=;�=��5�F�!,��xS<����fi��� ���ZJ��%��C���iYx���R��d��C����3x��a���/��,��:�0��~���D[�Xט��l���DB��ZC�N��(�!$C�������N�x%�aB,���ݷHm��4�sƏ$�^��=9�P8"��r��n�T�ǬO�����˄)s]�ǿ��Aaw�;dGò�q���̠�`�>2ǆe;z�şqS�yX��/a��
d��x\�PBB�g�z�Y����k]� .��I~?T����j��6����Y�k���bL��=�I��f1�� ��h����v�m� ���E7�?���񇷮k6~����T��l���F��E!��l�Q��~ ��	���y^P5�Z)�?d���7H�كr���R?z�2:9
Yo2&n��9����̡����6��v~��������+�]�_�j*�>Ix��:�N�uՈ=�GK$Ա�ec�#N���������}Q�����f�9NJK�d��R\Z��1hA��)���C�Pr���p����'v��.MW8�"f�f�Xhc�_������o��5EJح���#��D9� �%�^ď�ȱ3�ܩr��o���D��HIi��D(���#k!&x�f�C\�zg���N'���9����\��:7����:	���~���Y��� 2p��%&�-�[C�!�c�Z*����Xo���z�p ����UŇ%Zo����_= �P�P�w���>��?K	W���0#�,�������9a���v�:\�s��M��?~a��W��񢓜��4��Ƶ��+�5�4����-��r������j	G���弜<���Ս��Q�����i:nO�_~e��]��z��EŔã%���XL��D�~w���խ뚍o�U�ln
K����L[US�BH��0_���#@��Ek��_��ܤy��vB�z��s2f\���a�G0&���������nX|[�-R�:m{u_�ʓ`ҌI2ĂrI3&�w:�^};�b�`��u���Ч8s?�2��Å�!n���Tv�\*��J��(��\Q-q| �М,�q,��q7t}�:�g�ƏG�Z��S�ں~�w�04'ځ�����h�$���87��קt��z���Ei�x.�*����HiQ��A_��W���uV��ij��ˈ1Cc��jF�����KW�>?y����������<�hDD�U�!� �y�a�߿wt-}х�ĺf���Y���E�pS���BrX>�Z��C��MU�4�D"���c�%%�3�� �J`Ʉ��dV�l���.}P[������eV��K˦_���3kL$��Y����eW���09�v�vq|�L[�2C����u=
��?5�(�	�ڰvM���>!��YJZ`=�����8f����Ht�:��,������];wXX�̥=r���>%��Vc�� %eu���%��J���:/nw 
� ��6=-~t[�tX�vu��� �%2����e%���'r��{2f�L)-���s.��&���z]�M��ܮ�G��}Њ��a����~<�O)A%�	
�DD��:�\&?{� ��c��Z*}����Gb�Dq|v�y��n��S�����U��Bf�=ރemH���ǃ�f���\�'��;���^���k*,}ϼ��%&F��^N��\m;穨õĒJVJ?x��7���w~<�D]W_ty�NaW��憈��vu����Ee���)� ���RZ1�vQ9s�}1j�T׌�&�*��ٗ������aV�@�`�	Q��������@�ud��y�$ی���I;��~�m�|rV�� 8ஸb�a�@[oͥ���J��5?����4h��cC�S�o�|cH�����C|���a�������hF�ˏ�O�O��i��8��c�z}N8fm13����Y*��"�������S�9(��~¨��<�o�z8��GyE��Ec���7��z�������9X�𛇤)^�aF%�еu�Q	�b�<�u���)u����	%�Y �t����}i�,���>Ǡ��.f[\Z/&�(gO�+-����q�IIi�tv�I_o����O�{�;�P�N !X���R��6�[�E�%�w,�ﺯtY�������/���1�|�d�8��+%��g���h^���&Xo�R_���eþ�YdC|Zף��P뿶���X�;�h���|���}��e��rN�DKK���뤭�tuu��+��	1)���~�QY��{q�b�3ǔ[K����=�n�d����ƚ�p�7L�:B�1�J��hA��a�L�aW��i�I�)9{� �?���Ĥ��Lm���Duo���t0��|��d
��q�h=D�]�����,���'�7����\���J���f���땓�ޖ1c%ma��^�O��N��*ɬo�r�zEW_�A2��uͱ��׆B᧜~���Br<�D�8��/�K
���?�}� �1�k����늴�����΁���W!�d7(y0i�͆���!����}g�Y��j�n�����y�����$va:6�R`�\�5�x�d�b�|&�.���]�#[�8��Q�BH�J��A�Y�d��(k�����3Ӡ�mEu����D RT*�+a!���\}�n���Ⅳ�且�����y-;U��lvMkHX|\ǉ�"� ��	�w�E%{h��uu��#�GOo5�����E3�v��B��/���4�όk(!�"5#o����?_^Q+�ܤ^_�xH�B�bє����&�ıX1ǉ��.l��x�D%�%􆣍��0E!��*e�R4�'�)�47A�-}R:bp����}�iU���"Ο�Z���޾��K�IiɈ���KH1~D!�xO8ҟ�S'�rC�!ގv\��{;������W1N*�[%U ��bib*Fn����.�4������e0R&&M�E��A�#[�8q���#�"_�����@!����<2^��¡6	������{]�]�>k�+cw�;Kef�j<;�`]s��k���@e���'%b1�'��fH�Ius�:B!�B򈯿|ɲ搐�D��&�2 4Cu�B!��D:��$%B���Vq�ِ��B4u�B)h��A-��t�*�: N�?��APZq;�����7��/a=K�Rݞ��B!$�h�u�O�!�xE!������ 0�wm�z	���m��zw?kmB�(q����뺯_HrT��E�%.�[^~K�;BH�PY$��%�2`���⠬+E!���+��$��M ܏^��jj��B�B�@QG!�� D���\u8vZ蜃~C��pi�	!����e��.�yN���#�B���X &�MkP�ސ�F�`��N�BH��T@BH:ٜ��BI���ar�DX0��K&�7���z�1�-�N\�F���_8P~S���y���:�E!�Y9�^�\����*i�*�X46d۪X�TI���B!i��	�c�U�u��]v[�t<�NTq�Lԩ��-R��6x��<�|�?�bжX���2-�}�D��|�D�R��`u���ie��:X"�Ȑ �*z�X?����^aB�VB"�U�l^���u;%(��F!�<t7����?\U"�G̒v	K~�F�TɌ�1R_\麝�!�||����Q�Q'Y�tH�a�v�?�g`�N��6�_��Ab�襖�k���w�L&,B}fp8_d}����j>?��ZQI�!$�	ǔ��
Qg���u�B����zۥ�r"1�®��V*J�=�w.�|��oӇ��a�J5a����2�-|m��ji��e{~a��c�����8&}�Zܚ+��gt_�<�4>�ϛE1!�d���S�f󴮭�f�8��on�����(�!�$'�������#RV^#c'��zWϼ!��.] `�3��Q�d	S v��Ѯ��7�����.��l-`~bv�8��� ���A3Ě>��%���f�����[r;E!$�)���$��uk6ׅB�-n>JQG!FOz�3��A:6
�[�����R�/]0d��P8"��r��n�T�����;}|�L�2��>{{Z%WЖ2;+�ov�.a�]�p�2� �jVЦ��m���ǂq�q��h���$��S���猯#�d+��ܝ�غ���F7V:@QG!Y&�:)��pC$������%C✴�&�n]Ոk��r���#F� }gʥ�K���ϘE�-�t���D��oZ}���k�������D�K��)�N[��p�i~㒢��̈́%�X���W��n_��BL�n���S�BH�0����DJ���D�v�3'��d[�@���;SΝ: ��V��K��~���VKQQ�J���k���H�0�3K&b��2M]EY�u���a�� ڍ�B� KYQ_�Q�l^([�5�&J��F�i@QG!Y,m���n�=�o�*�ރ��v�H�O��P("�&͓����sU�Z�ɘqU�%�I>��tN�g�GB�}B!��&nj	@�A�E�Mn�.5u���������b��=�o�j�I$����Hoo��DJ%_��Ji�V�T����%����K�ߖ1�u�l��X���H!f���}ts�_��p���.]A(�!$�Ѯ�p��r�gd+�q�DN�|Oƌ�)��5����t ��M%�p�L[gFתõ�u��@G��g�A'OA;*qO�̖�w��#��v��U�����'��*+�-k6�$EqCg���B����zx���Kx��02)e��%�Ҋ�2aRHN�x_F��&�5c%��צpis�:'�"��ە��>�(��|LUV7[�(�]wO�ډ6���LQG�5`E�b�k�o]��nl�޺�t���Ѕ���*BQG!Y&��7!6�Ƅ>�K�F�"ŵ2a�r����r���w���VJgG�tw�KG�e�]o��I52���޽�u�g��u�F�$ ^,RwH�)�%ږɲMHv��e��Ue'k���k��5�d+n��$Y��쌦*+��dU^'��b{[2�SQI3�K6%Q )RE��w�{�y�n6�@_��sN��S�>�o������v��t%@��_n��Bz����������ņP�3}O����oeQz�~�:m[�����p��4 H*mw�l����ϳ������ηӦ�MM;r�pW�a�#�@L�~�P�͚e�=��/���
j��*��knYk]�A;3zԎ}��M�6?7c�T�֭=;�j6�T�ۛ�7�W>��t�s���_�|~ۊBzl���O�*��a,������������i�80�ʫ��7_�$S�KYz{g�=�U��ڀ�2������6m˅�n�Z��q�����P 1����j����cbjɕ,} �֨��W�Tȋb�3�����2�5;=b�G�"*g�K��c��t�c�!�/�R��r�M�����3�v���3Xd�R��9���{ k�ͫ��G����v�s/�Q��1 �$.����v�]��j�'�P 1��AA�����2����{����w#w�(��uZ��y����}MXSs��F�g�֙Ry����
��z������n��_8S!����\�.u�
�? �vu cj$�\s��qK��5��2����q�W���*��ī�L|U�������ﱗ  A"�@���-5�MN=3>�ySKl_�˞��^w��0���vk[�9����옵57Ys.�Ukzn���3�n�bm��/����{�  @eu s
n~�O8pxq��V\jޗ.��0�����/�~a   �u �R�p�W��+)e�  H>B    $�    �P    	F�   �k޴iӖU�VE� Z[[������է��   ���:    H0B    $�    �P    	F�   �#�   @��     ��ޛ���eT ���徎[��Z�j��ի;g3Y����c�T}�Sٴ�6Fg�   �W���s�����z�W֯_����ı�U�����7    ���K    H0B��L��`G�}�   B��d�[m�k�   <�:    H0B    $�    �P    Q.;��u��~�����vz�Ł��   @b(�m<9hI���ӹo	,��    �Ԯ;>d��ٺ�졲nW��2��    Ԍt媧@��u    B׵�����{��6p��\sYɷ��@��u    B��w��Ĕ���?Y��?]���9�y�;B   ���?���~���\t���t���L��m|�ƲoK�+AKK��}�n    *Rn��5g�������r�5�<��/�ۋ߷q�   @��J������7t��w?��^�2    ��k[/��_eMM����Դ���q{湷,w�m���\����N���=j�<��B�+����a�    >2Y�3���eK����q�'��С���_�;?og�L���P��׏Y63oa"�   �;~|��o�tA��+��L&��)�P�?>d�ׯY��#�r�6B   �:���ǎ��|��K3��w��(7�@'�:    H0B   ���}�G���     �u    ��ɡI���;粖t�Z[[�-��H���s�mj	�\!�   �o�k�O�wy:�d]Е�)�����;�r��(7�+w���P    �R�-�$���c����l�K�����fs�Y׺�&B   �D;�����7;r4�r��x䰅�P    	F�   �#�   @��    ����]ikϜ�F�I7���+�-�   @,��pq��[������)нv�'m������    �V��j��    �Z�� ��    �^�����    $B�� ��    $�v��;hIu��P    Q֍��Փ#�TkΜ���:    �C��Ɠ��dg��޲��X=B   �D��@��u    b���T�#�   ��zt^��P    ��9�y�;B   �X���+u�<��֏��ڍeߖP    �֜�F�>>L�   �FC�   �h���B�~�U��T<�LMM�˯�g�{+��"�   H�L����m��e���G��i;t�e��(��   @����ö~C����Q��z�2�L�0�UT��
�   @����c�mn>s��+�r�"�   @��     �u    �`�:    u��ФM�̝sYK:c��-uY��    ԅ7ߵ�'�λ<�n��.���N���\�P    �R�-�$���c'���3�pU��u    ����K8j���Ѻ(��    �P    4{��zo���V���������d�   @(�~�N�'����OX��N�uǇ\����'� �   �����^��G�x��{?�.Wo���rN��J[{�5�L��F�_X�m	u    �s�e[z
q
y�.��]���sz�Źo��z�@���������nO�   P3�C�e_����@'�:    �V��.�@'�:    �Wo�.�@'�:    ����a;n����/u�8���)��tB�   �SW��Z%���S6�wВ��
,�	�   @�/�ޟ���oS�uc'����w~i�/�@`�G�   ��S#n/��]v�9�xrВL���Վ]|} �G�   �������ꮅ��!�   M��6���	�z��e���z���-�����+Υ��@�]�喪��   @(�]r����.�i�q�t�����l�(:��D�#�   E��?�kn��+�]w|�:��)�)�����N�niPρΫ6��    N{�uo�t�.�����w]�{�����i�{��W�>�y
v3���˾-�   @���J��y��PKm]���^���U��ǚ3C�H�Ǉ	u    ����׏�C�   ��)�]C0����)�g���۔�׶^h�o�ʚ��Ǜ��i{�����soYP�*��   @�|o�F���'��K�7����[�ߦ\��ٙ�Q۲��Z[Ϗ8��v��Q�f����-D�   8��i>���-��i�KͱSo���=z�����ö~C����Q��z�2�L�0�UT��
�   @(v}�	�3�P��
���_8����r�x��*���ǎ��|��K3WT�E�   ��6W��}�G.�:�:    �Q��6��(�s�4�N�/�KW��8JG�   
ma�M�5gN
C�.�1����U9��q�    �B�(��!�O<{�������1���){��̓C�6=3w�e-錵��X��*Wu    �a��[i]�վjq(f5��1��?1t���t�]tAW�pVT�z�:    ���2�ݯv�-��B]�6����e�+�d��؉a��6\EUn!B   ��OL�x��=�Ɓ7��pԼّ����-D�   8�4�n�P�B*�@��P    p~�V�\)��a����    N�ϕS�R���חB`5��42B   �P���nh��,����F�u�:��~xf�x��]�!�Z:3o�n�m������nK�   ���i����;o�7n]f�i�����-4��n�]�ɺv
t���oO�   �5�S�/�3'
t�̡��`Wm�B   ��P��d1�zvA:!�   \����K5p���0�ނ]P�Nu    �@���O�u��G�V�,�^�]��Nu    �a�Ŷ1X�6+�����;�T��rY�   @��G	��]��(�u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#ԡ*�O��G^6ki���dldU����   ��UI��ܻGlÆW�m3#�  ��P�3gθ�qv
t'O�4�p�   ��P�@�`���iq155e�N�2   ����������1   ���-����Ӂ�_{[��tz�   ����6������V�ܴi��ޓo   5B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�5���_e���N	�~���O��mz�k;3d  ԃ�-[mt�U��:4�������\`��~z� �����w �z0ٵŒ�P��06l��S��x   �"�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:4��-i�⥭��ߦ�������   Q#ԡ!��ͮ\���6�m3    u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P��0�1;8�	��F�L   �:4�S��Gf���#�   �:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P����)e���~��Ρ   �F�k�;8>k#��@���l���u�)�� CݦM�u   �B]�8xf���ա������   ���     �u    �`�:    H0B    $�    �P�Ě�����)�d2���d�W��T*e   @#!�!�����,�ͺ���͹�u���   �PuH$���@�)����X[[�   ��P�DҐ�r.   ����9tn���   @#!�!��(����9=s---���j   @#!�!��JGG��C�W�$�  ��X
v�.�rl:c���Tp�x�   �8 �   @�����q;u��Ess�uvv   P�u��ɓ'-n�w݆   �W�:T-��N�����v   P�u��l{��u]`]�.���fl�}�   ��P���n����{-�f   �O�:    H0B    $�    �P ��ؖ�6ٵ�  ��]�-Iu ���n��  @4u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u "u���?�j��Z�lr|���W߱7G��> h<�: �Z�����T��e��Ykon2��� ���     �u    �`�: ei��#G��d0�FO���>bsss��MNN��![31S��gfglv������X�>/~�)����N<�b���-��,^�������W}��S�vf����}� �x��Pw��w���ޠ�o~���-W�u��kÀz� r�/���)[7L��>d�����uZ0�^{��_�/'���P}ڤ����]�7��`J�3��5{��]} Ш�6��(��yPw�>i-��r�PO��T ���ٮ��zkoow��袋������>|������CCCv��	�Fww�vs1
"���U�V���DC�'  ���Cݢ�����3��9rĀzSm Q������mݺ�.��[�~��.�`���y�fggmffƅ�~<x�~��_�L�D�P�
z���� ��5D�kii�իW��U@�K��O~�~�7~�� �.?p^SS��]�v���7o��o���8���ةS���^������z���� ��T(Lz}  c��0���G��m����*i浸��[յa��f�-�И��o��� r�ڗ��%��C���J��
&�y�ץ�^���v�m�ٱc�\X�>�"�'  �.D�Sǭ�����!YRss6;9i-s��8;H�:�� 
����k��~���f��׍��K�N
%���'���_1�DD*��/��.dEY���/�b������v  D�!B��h.I����5kָOÑ,����u۸q�ǩq>::z�r���� �s����	s��%�Vٴi���SQQ )��A$���!�q�O  p��ujt��4Tjݺu�a�dч jH��4I��S�+5�h�������=DԋT��QHa��+�t���ۿm===���]�A�����W���Q�  �T� ��� ��G�Gv�w�@�!���\�e~��_�����+��f�>	v  ���Sj ��+�����2�q���Y��'O�^�k���y�%�#�P�;  j�P�� �}�v��?����I�ya�@��O�ľ��o-nĝ/� B}�  �%B��J w�y��ܹӭ��\�ri��B���z���/�2� B}�
� �� ��� �T~я��D�O�  Q ԅH��k�˹��Z��A>33��V:.��}�)�xa�` @Tu!v�;��K�m���J���_C{��뮳���߯� ���g��7���q���l}>���gϞ%�#� BЀJ	 ڣOa���'n��JD.��"������kK�A$���e~���?��l};v,��  �!�huk��72\�z�n�!�Z�p~~�������̙3v�7ح��jO=�Ԓ�)�=�βo������p� �  ���� ���O�n��7���w��7ߴ���߱�^zi��`Ah��ܼy��a�'  8��9���j�җ�T�D4gR�n��u�h�����K���_�> ��u 577�=����!��a���\5,R��������4b}j~]X�	  �F����o��۷�U=�����p�|�w�}��/�l} ���B��H���h_�z[�g����`����~Gջ444d���'�����>��`�  G�Q*�r�h�m.����s�aU?�2/#�%׶m��p�F�U�BN�<iw�uW !���> @q��)���<�b�I�Z[[]��sW��A��g?�ن�U�|����ȲK���> ��u����][[���k�mRhԍ7���A|Æ�����>���B�yVP�	  �G�C(ԛ711�z����d��$���>g---�Un#�.��N�8Q��P�gU�  `y�:�J�0���\��B^�a���f����:;;�رcv�m�������oO}����  +#ԡ&�&''�'��wG�7>4�Id7��Գt���馛*
!�繪�O  �2BjJ+�jHZ{{;[#���?�qzO�h��ߐ\�nccceݞ�<W��	  VF�C�)ȍ����իݰL���*��_~9�A���ڒ����%ߎ�\��S�`�[�  �4�:DF�1�"*Iok����>粗�o��Sc����!�R�h��+�����Q�竴> @iu����t];=���!K���.���K��U@�e�֭eݎ�\Z��	  JC�C��%�%х^ȼ�"�������,���  �!�!���Ӗ4�k�R�>hа�rP��UR�  �4�:Ć��iULŵ���|�Y�����Y\%�	  JC�C��`�>v��J��i?E���y`�<�zI��>���> @iu���MMM��Q6�������cY���  �(�;�ӧ��   ���f�繯�l:�|�l8��tֺS��6�ZO*e7��Xu�%��i��   q���e����_�v�u�kj�M���Rf���u�%K  @\(�ͧ2{��=P����3ۛ�i���r�.�'�pG�Cli^�u �ѿ��oڗn�΀ �N��]����K�޳��\G�?Ͼf��OJ:6k6�ͦ��=���A��z�v���hv�n��P��Ro���K������d&>���ˇ��o���^��9��V��7�x���P��UR���/��8�\��cU����>�����Ѩ�:bK���������e��5E_�k��N|c��>�}��s������7��t���Y�]�kZ4%�NǾ��Ԧʟ�;���[�Z�9sư4�k��r��,����W/ƨ�GaN��8�\G��t~*Ѝ�gz�����3�ܽ������Lz��`G�C��f�<�B3�7==]��N곸J�^��3���3���6�����M��\G\�t����7�^�����<��u@v��s�}��������nG}.����gjL,נ ��:�Fs��3;j�<�����6Y�{������!�I�r��	ۼy��W&'�·<p�@Y��>�Vi} Pk��N��=X�r5���}�*]<�P��S��*����������]x��o���q[�v����Keݎ�\Z��	 @-iۂ3��U��s�=���J�a���_��(�h�JB�+��B}��>�ֽ��z�����z�  �mz>��ط{8{_߮T*�p�7%�!���g�yƾ�P��3��~��n���O�W��U�sA��5��_��^?b��F P��Y�~�.i�����-���P4��'O��N�^{-�挎��ᾕ��Ҽ:��W��O  j!���[|�[�s�uH���GC�^x�����mnn����uvv�O�ӊnO}�����U�g\t�nsC1�����,#�������.y��^�]�}��s��]w��n+�ձ�Cs���y�}�C�.`�����/9��W����7]m�_�t�Ǽ�g�������=N�I�<��	C|���?�W�����λ^��^瞽���Z��v���%o���}��ӹ�O�n�ۭ�^Uʹ^x��K.X�L���'�]�,=Ϟk.[|.�>� h�K-Tb11����d҄:�z<���O�=����C��z��ۦpV)��,էzYM}����h5h�&9���^�2�0G��>�#�X�ԈU S��u�.�u
{���Fr�S����]c���j��q�k�z
t����K)<N���+�qc��x�y�����U.�K.��^�R�\ra1wN(�W�*�\�?�{C�;�����������_�^�<��dm�bD[tܿo��!��:$�B]SS���������SO�G?�ц����{ϭ���c��1�>�
�>�QC�	O�#5
{C����rz��^G5Luu-�֩q�Fna#S�X5�ըu�s`}w��5�������!�u��U#</�U��u����a�ნ�PJ=�K�:��
G
T{K8G|��,(����s]���u|�{�������?�=��\�9^��J����ō�f��.�pB 7L�?��m߾�aC����
j�o��4�����>��8���,��@԰�A�5J�xv��\#:���5t��o��P���hw=u�������{
���!��{������F��:��Jy�ѹ��T������[ι�WK=�bCKWR��J&���Q�L� �뗿��k|_w�u9�Q�h�����'�ܟ�S+a~��l�`t}�� ���z;Dp��z�
�\���?�R��+�=�Oe��}T���^��R����+�Z)������T�ܳe�#�uC�B��YN�+�\_�ia�f���"�!47�yuᚚ����뿶����j��`
]
!���r��Ͽ����o���L05X\/�Ĕ���G
����<�K_5�ESw�BC�ͽ\��+��a����\,u�_���{�D��`ņ�\԰��#����W˝����A��z�^a-@���_%��������T�a��^��:$F�0C���7�\�cǎ��ի]�l}.E_�;�F@>�*�]�5���䵜��`.�R��0�{���?S�<*}/��Q�B)~�}���'&c�=j��?7x�綐��/~8b!�G�78/���,�}��s��{b��K}h�ܪ��Y�y�|�:$��Ԇ�=��Cn��64D�VgԊ�~�i���p�ҩ񪆈�����_V������]_t�g�B:�PWw�9��ł�B���o��C�<݇�~5� �I�~�(�����z+_Ƙ�S������9���ߋ
���M�u����,�}��s]��yr^h��w��4۶q��
��L��ҥO�C"dzY3�N���~���.�s=ӰH�T�����|'�2���}�j��3�O�Y��q(��!
{'\p�}�o ~�\a�ׇ8?�-(n��>�zF�CS��<��{����o���r�l���m1p����Ntn�+<�6�z �R��{Ҋ�GW���BŞ7�G�C"�|��Z���/�l�z�c��������v(��y�'�\jh�p���r�����]�6�2���0�{����[e�Rz�s�@��o���Ph�[f�e:�ԳV���Gt[d,(�Gn�\�/��R��r=���=��7�x��n�VU�g��J,����z�b�S�k�n+�xB��g����v��׻/4���l۶�n��&knn}�`~}����e�]-�s�̅�rC�)֐J��]��g>rvq;��T#x��N��a�����Vl��R�p�մ^�7cY>�-L�������W��=`~%�b���=�Z�d��]de�����:��A��Be�|b�g��C��&R�S��:Ğz�OW{��1��G>bO>�d]���n���m����裏֤L_�����π�O�}�F5DԘ��c���QH�G�׿U�m����_��b��󸫄�I�W��`�J!;.d�PJ�큘w���JC6�r��r��W:��y���CQf�
[�}�R+k�BbO��h�	ԞBH{{�}�pAdvv֒n˖-��/~������d�W>�gkk+�����n��S�������\ H��Y����v�����͙toٷ1 �O--|�y����$���^��K\ �bޗ�^R�ɡpX����߽��}-^6T?=� Ј�Y�b�rz˽��F���zvq
 �gr��'BZ�+S�����F5�,�@�(@�rMλ�v�uO��=��Xw__�z˽���E���]j�߻��VOD���'>���	�"��[�e_|ql��s�ƍ��O=���q���X�ƽ��Wc��l�<-��a���G��޾�D(A+�2�G[S��"�_���+�J�䦄:�ZRz����;���-[��U�V��>�1{���ȑ�/@���cw�q�e2���8�P̵k�&�>{,���4�o���t�?�-�}��{r{2��~�o���
wn�gd	�V��w����Ҿ\Z������(@�䚝ۣ�[�ќ�SI/��[---,�CSSSv��	��[\O�+����Ԯ�.�o��W_mo���=���G�@`bb���F}�G�c
U��������Es���[�ma_1��-?�k��ƾ.c	�`(4��L�ڤya�������j����L �t�}=���|-�U�����ޞP��R/�z?z]�p�M�6�s�=���n��Vף������~x�������g�*]F��Q��ˆkX��zs|O��S�SO!�0�燺��%�wA:���{�O�)k�O��ξ۷{�ej�t&Wfu�%ͥ��.���v:�v~��2��)*�/M��뮳W_}�~�X�P��P���!s�s��
r^��'  ��J�MM��;��Lz��a�����g���5������.G�S��52�k�f��뮻���_��4��𡡁'O��|��jP��ѐ9�ysA��#�����E.*�6�^X8C�mǍ[�����Ш�4Գ��;�r	� ,����k(��\����@'�:Ďz*��hs��to���<x�:::�s����Y��)Z���k�uy_q�v��i������˙���t��o��g�J��Ri(���K�+ĉ������^5C45oם7�ysn���B
Q
z�c�r�������������=��
7|�ֆ�Q�	 ��ԋ��o�{�k�J���}]��T<�����@e]�ɤlUkk(C\F�x�7'��nsaGC�4G��@��^�_��_wD���>��[92,����z�5�\Mժ>����ի]��^�T
X��la��k��G=X�S ��_E����_��S�{�����O.D�Ebr�ٯƩ���R�/%�ߣ(@2�-���uܷo�|*�g�����?�]���-@�:Ć��Ԟo�;�����W��Ұ��f�n^�(�|�����v�����GV�_j�G���/mr��".��R�k��"r~��[����܇ͷ|f��jU����YAY��~�z{��W���{,��Jܐȼ��n�d�2}�}�G�-Z�zs���_�>�|��[~/�׿��u�.��Pņ�Qn2�V���GV<N�r��@mh��fK�,�~��L�ؼ�/u��65omjڑ���s��2��������+��ȻvIg�FFFB_eT��رc��W������W����y�fף��ﭷ޲�G���ZR@�ܶuw�w6�~Ӳ�FU��N�էz�4�qfff񶱨϶ա��`T�S���D���W���PV��^{>��Bd�P@?ɣ׵�zM��<��p�����f{8����Ke3)�?.�mږqݖ������q��S����5���[��.����̴k��z	8�t��o�iq�zP������ r�m%����e���LOQ�*��j9�M�N=cjt����]_�=?|r�gG�R�S�~ΠGa�R���zE�U��e���LK� z.����v�]���RB"G����+>�ֽ��5�N�BH�-�QK�]k쿽�s��|�O��읉�����1k7�\�QK]vm��\}��U[��P/�B��WM
�P��ڹu�婜Z���Q���ϸ�Q�79wC.s�_ϱ^�Q�\ũ�L����~�?�"B"U/�Ns�^��K*�J�%�쳿y�9�Gh����e�Ƈj���7r7�炀��X���9�[,��E��nS�\��:\=���.|�Q�\ť�LHh�U�s � h�:DBaNC�V�.)���ؚ�v���� C�R����q,�H=�@�a���F�蹪u�~S?S��T�z���:�\nOI��M��{T{[���,ן_���'�5���^˿hL�C���{����#�F�_�R�/saÅ���!U���蹪u�~���v�EE>�y�|���U8�Y�Q����>���^g�ޤ�ʿ?��ms����x$��+}H�r�3��C�׊�"�HB��E��n�΅�W�{��&�b뙨�P3������ ����O��x^�����M̱�E%�>����C�G<���yznK��(k�)��TY*[�}�a�FLX�*DUn=WQ�����ܗ�p��^y�� TaG�K�g�;{�x��:�s����"��Q�QL�!^�W8��-�p476��k�Ø��-�*��q��u}������[����.W���?��~��^ޏ��?�A�;���zE�CM�;�b@�����`4Z}��Cr&5��/����	�f�¥6����h�o��j�y5Pܢ(���k�}�3�1)Ć��e�Q�\E�[�yQ�CZ���X��X�7nue�įt6^<o�ӽ�_�p�[�=e>䨞}o���?�¨g=W����P���|���*pz��<��P�P)�i�z�; >�'����y=F>�(x�J�qmp�aFn��\�M��Ay=�E�U#��E)���qs������~��^�b������\����z��ʵaЇN�}�=��ĉ��> ���>�C�g��.Ե��~��-H4����|�P��)�i��0��"ņ �rטPO^�q5X��X�<�c&j��b�Y-ʍ"HG�]�7�WR/s��S�>ȅ߻�7M���6�p�@�>���d!�[������Hi��Fa���繑����U����;�T-������z,n���ߋz^��P����g�[�<9��0K��[�P�b���\j�q�O��	�c�a�]~�)z�~�q?R�*�O��*�P�v�Zͮe��R��z�%��7?�i�!�a.���O�]�y�����p�?����ͽo��^a���
�ş��{]&a���ɇ��^c?3L�����ܞ�C�5�U�ר�zF��z��k����)+��9���8 ��FB�m����U4&� �'��F�_|��SQ�l��A����Qܜ�\�8�����\X^���y.����De*$�h�����sɯX���lj��U*��9F��?o|�Q>/�`L�<�d�zN����}�E���s\�%�5����Ι���{~�d͞o�u!����Ş, @p�<�\�*�@��V3��7:����A�:��[���WI�����q�XT�_ �phg��}A�勢L)܇p�,��W��
{��X�)�*��u-,7��^��*W=Xz�U=�!��Baa��Z���3Y�����#�: @"�/*��e��s��~uK?���Z�����*2o-̍�����a�����'~�<?-��/k]��� �����
�;��!��N��[/�F����P H,���Х��9ao6��?�%5N\�]�5S ����Bm�a��i��ד��	�F�~��r=Vn�b�q(��H���|Q�%�K��É��n�\ʭ7>��gB  �
����Z7��Z��HX��}��6Ȁ�XX��-E�+��綰a�/�os&�x�S���(ʌj�Z�y�6�Ν_n���s-��E����r���P H$�s�����\�j����σ��\n�Ͻ��+��޲��\�
��_�����J��T�]����.���	jq�(�\NT���-�s�틋���R6�\ʍ[�Q*tB� $�r�D�f��ׅ�"���x��v���ܼ>y�߰��9Uf�\�P�ϛWX��w[F��s=�R��"4>H���'�Q�����!�_�ޯ,�K���:w)�r��R�Nu �D����Ԟ,~>��G�c�sH�z�
;~���h��}��\��y.X�\5�t�~��9�z˂|�(�P\��_E�m�P��ԝ�!��\ʭ�ߣb�Nu  Ĝ��V�e��>�x�r��;������[#���}��|(势O?�0_�\�$�)Q�?dY_~�B��~�iX[�P.�&�r�Nu!�>uڣ��6o�L]��OOO�xܺu묵��  ,n���?o�u7��,�^����-����(S#̇J�x�\�<�2��0.|�s�2���Z�F���+:!ԅh�@�����Y�k� �M����Q������Q�r�J�
�5쵪u���C�h�W��e��\ʍ�R��   Q5�)�r��@'�: !�Y�y�k�R��L��Kg���R���oO*e7   ��@'�: �\��L�ؼ�}���9t��ж�����iG.��J�]n   H�r��R��Oe��?�{���N��=8m�7���u����R�=�;  ���$�	����/�H6��3����qc�}�;�]��i@ >�y���͵س�Vʥ\ʭ�ܨ|�חr�ܰT�!B��А�>}�&e]u�U�?oܸ�ZZZܶH��A{{������Yss0�F٬�0ה�����-H�v���Z{�@����p�i@k�N����ǼW�}��C��K�+��܇>o�����[�Q�U�!B]T�����.yִ��ի�=nvv�2�L��)Ѝ�gz��e��U��7w�o���9� �  �C��Nu!���6�z��������B�̴��^�e���u����|��^���H�  �� ��6B��ު��A��C�͡Ӑ�0{�
)ح�������3   D"�@'�VBD%c!̡+��bvܿo���b�!�AI�Rn�1�R.�_nT2���[G�!�@'�v�m[p�����*t.���9��0L�D�Kgf�mbb�����͛��ň(�r)7�r������:*7hA:��Pw�С�ܷTP������fK�̀�L�gz#} �vg��ەJ�6`�$���٭[�R�T+Ɩ�G�r)�r�/7*)^_ʭ�r�F���u@�e��}m���>v���KoJQ���?��K��[�r����K�uTn��
t��w��dR�~��~cnJT�� ��R.�Rn�����K�uTn��t��w ��*���Kg�[2iBJ�?�'O�����ߺ��@��R.�Rnr�mM���[G�+�@'�}w �*k#Z}���}#�D9���sDK�t4��
�K���\S���[G喪�Nu@�e�V�-V�����   ��U�BPc�tf�bFA3E�  D-��      �tB�jl|.~�/�{����   *E�B     �@'�:���4۶q��
��L���  �"�   @��s�b1�K�l�   �u@��2@���   �H�:��b���ۖ�X�e���U�V�t�5k(�r)7F�F��חr�ܸ!�5�2�\{ߎ3�ܽ�b�9��5���x��u���i�\ʥ܈ˍ�^_ʭ�r�PD �uA*�.�׀���͛˾][[��^�Rʥ\ʭ�ܨ�����:*7�u@R)��mg_���݃Q>�u�����ЀT�ԫ�)�R.�V_nT���Rn�g�: "mM��i�p~�ξ�T*�׀�R����z����P.�Rn��F%��K�uTnꀈ�ޗ�G9���9��^:�"�N[ss��:u�r)�rVnTҼ��[G�&��P������L|c��,Wa2�vP�l6k333�K����r������:*7	u@��S�<�}=�o�p-���L�L   �B�T�n�hJ�� �)�5g��  ��: |��{��7���r�:  @}!�1�`�^�u�}k�؃_nUʝ}]��0�+:�n�=���/{̧:˟�>4�bώwX5(�r)��r����~�ߣ��Q/Z*���oߎ�Tf��7wTsn��t���H��K�	-7*���K�uTn��v͖�Y.��<k���y�_�|;mj��Դ#w�   ���1�����w6��Y��X*3�I�`�q�lӶ\�붬�h��~   @c �	�^���nwޕ!.e   h0��inS���    
e����&ԕ!�B�pvh    �IY(�R��PW����S��3    �3���GU6��c����}�y3    GC/'�����Dط{8�{��T���     G�GY>��Lc};�hch��   Ț�Ӣ�Q>B]F�3=M��   иr���o���� �Ub���ѝ}
v���   ����.�Nu�R�3�Yw߷v�RYO   @.���Lo�C.��4�����ξ�uM�#e���   P?�r�2��曻�[���kQ�f핹    IEND�B`�PK
     `_[$7h�!  �!  /   images/a7fde0f7-2836-4f0c-aad0-66dcccec46ff.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     `_[wJ���  ��  /   images/f9728bc6-2422-4ead-9082-90351081a874.png�PNG

   IHDR  �  �   )��   	pHYs     ��  �8IDATx���	��e}�����sN�{���  �NpILbL&���'&HLn�F�u��%��Y43sI�b���q>���I"��+��4�4��Yj뽧P�j �s����?�.h�p��_=���   8�:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @: <�6��䪹��|X�&�L.,�t~'M���L���t2�ٙ4�	�l6M�����l(uBZ�>���f��?�[NL�~2���o'� �d��L�L;�]I�<�o��;����W5 �: <��û�;>-d�K;�lX�f:K�>f'�t8��p;mW&2�b�s(>�F���7|⍍�dj���̤���X����ه�$ݒ��9�z�}���[ ��@``�n�f8��8��ɞ��U�L�|�W�E�К?j#�2O�7x��I�B.������?|V(=�p2�9����O\2��d���Ω�8�J��d�w>o�����F  9��@����[.��j�ON�:�d�x��Ei��B��4�	��!�6�������k�ۍ������U�|'w&��]��Z|u�We�� `�t ���^qB�&���3[��QI6YR�4���1�b��<�ւv.,h�p��z�D�ُg�o�إ�Z��s��ұ��^��� `�t zڍ7�X�w��gwBxq���ʵ�ݛ;$���I'�)7C�P
ݏ�������o�̵��϶r_�w�m�λm���I  
�@O��o(ݿ{�w�'���;�w�|b:ӫ�I�ۅ�Px|��5�ڹ��'��\��F�������� Ϟ@ z�7zd:+���֋�Ӹ��d�S
r�l����Cn�^5��?ټ��$��N���w���� �� Dg�������$���������ڒ4�D03������6NitW���u��Kv����3�]5��nZ< <=�@6|r�±�ɋ���/?�}��N�Ƕ����~|�\�!�^����_\�y�w
��?e�e�n����  ���!s����/,��]H~��c�v*Β��N�S�����\��͗|���ڕ��ض�n��� A�0�F7]3��=����B��zh����N>�7�W��>f��K6��F����P�|���� (���ۼys��/�v��^=��rb'c���N�^��
�l�����+���r�k6�S �#��6����c�C�?���g^���&�i=��X??��o�؟�e�U�����߾��Wo 0 : Uw����W^��4.j���f6�3�ʶ�J�ՙ��W���5�*��[FVW>zU�N �>%�8(ֿ���uJ�?�T�3��ζg8���5
�S���'�oY����'7��o_���  }F��ߴ�7ZC�׍g��2�]�L�v�=��]U_�}�%���Ul�޵񢍟	 �': �Xw��/^�(7���luE��]U���¦7}������{g����m��	t ؆��0���n��U�B{~�C��k�l�64>��㵷���\k�/�ܽ� �$���4�w�G&�ӵ�w��;i;@dZ��⩏���^�=�Z�_���� �C: O�M����K6^�]��V rIhM�گ��/[��u�+����Ƌ7> �t ��+n�bE����z���f������d:�j���L!�+k>��S�f�τ: ���y�Mo=�Z�_1V�xY7p��4����K����~h��.7����{��  � �7�����{J�^��N)@��d;��R��R㗧B�$�����k�=  "`��n�f�]�q���دw�9��J�T]�[���������y׬^�:	 �0��}`��kC[״Bkn��d���r�����k�?��~o�� b`��}��_h����Dn� ��m-m�n]{�G.}�Hk�������z �CD��� �ɡ�_W���i�	������5��O�ټ����ٗ]��v �a�����7�����?�3�o���� <�4tr�B�ōv붵������v>��$����M���=����j��I2��r�u�%�������k��� ���n]�*&�O�'�Oӎ���,�r�Ò��Mk>������o����  �H����t��Jc��
h;;<7��f���Ks�>���ѿ��5? `�t�>q�M��i_?��<9 U�K�Vgծ��Cks�МK�`:t��!ݐ�����R�u�L��i�=.R+�/h�[�^w�e�_w�;�> �A$�zؕ�\y�O���z�~x fD;�OO��K?��?d�7\���� pt����+�x_q|m'�)xf��䖍,���M���$I��^p j�ک��ֿ��e�o��h�� �#��c6|r�½��7���� h&��I�O,OUyw�:٘���KvW��w�v'����b��O&	��H�/�l^����|�-��b�; Ϛ@�!k�7�k;�=�*��8H�Z:٬v��C�����FrݏsV�?��4;;'w�wN�l?2�h�ښ�~�{6�Z��x�Q�n[��+׹7�gK���7�wƯ���/O�Խ�t����U�U�'��B��]>kY��q����ڵ��M>�~trg��nX^��ʶ%Cc7]�������Y��\� ���� �]�=��Yh��˘鲧���j�����|%7��v?��ҽ��ɶ��[�Ƕ�j��@Gi'���P�5�G����׵�����o	 p�:@�W[?���`��n?˿43�2/��8y�I����㱾ml[s�16��^�7��-�r��+.�x�;�g � �"t�7�=瞿�(���-�̄��x��4:�\)�\�>ݳ��/:��Q��%�Ƿ7ܷu W֓L{dbx�������^���^ �g� ����+V|����7�ͣmig&��m/��􀶹���ٹ��ʉ�N(��j?��ֶ��[�=0_ٝ�f'K�՗|d�1Ci���^}��  OA�Dd���_2>T���m�0�v�v'S�~������-,t?N^zr���#���jv����m�|�$���o��[��o~�o� �It�H��������7v�L8vM>�s�,��g�׷u?&ɖ}[�y���Iߗz+�Z����[���u]��  ?ŋ@�Clt�5�����&�p��M�N�油�{0Rɝ�䔡���nݿ���]�5����N�S������?c��YW���'��������G�����KӴ���V���ys�|��yG���wD�{V�{��4����������b�U����Kn��w߽��c �@8d.��������i��ݓ{���'��Y����任�o{�oC�Ql�\8,�?/���W���Wo <�p�}��M���I%@DvW�����S��;{���'4&��v��xp��fw��ߴr�����y�6�f� M�̰�}C�R��08b4�Ix|1;��9���{N���=o��J��y_�}6;i�I;�̝�ݼ~��7_{�� X^̠K?��/'˓�H�~Z������ɜ�^#T�ܩ�N:nѱ�{����T�������Y���nY�꺋�{W ` E��/@�ڰyCqof콵|�� ��]�]�?��/?m�ǔ����C���B�HC'79�X��C돾���] 8Q���O��|�=�������s�G�;�"6\ɝu�Y�G�;���G�]�S����Ӵ��,U_�f�9sk���`�t�i��}k�Ndkk�G��"w ��_|����w<����j����#�G6l���V_� �0MF7�.�7?�ʶV�!�V-�6��Pq(z@�z�峖��ZZ����7���z����R�P?3�3��oX��W�4 }O�L����^jn���%zЮ�dUqUO�2!�9f�1���,/|�o�v����J��k��W��'G7]�/�|2 ��:�A����=�6���8_�G��i����zP%?�;oŹ#�M>ֺ��ժ�ɞ����5�O+�ӛ���W���޾; з:�A4z�[N���}0�&s�����=���xxq��������߷���^�?��o1>>1�i�U/��X �/	t��d��ѳ'��ޗd�� =n�1�i&�N1Wʆ���2'.>��b���W������g+��k�J+῿�����m�}�� @�� ��^q�D���~���7Y:kiO�f�f�^|�G�C���w꽺���7����e�/{�;W�� @_� ���������ć�L{v�>����=��'�"��������}=Y�\kI5>���7���?�jO �ot�����\U�5y�T��	��/e�F�{������.�ν���ܳ�������H���r�^߸k�ޏ�n��妻���,u�9�W7�2�a �2ݳ�'���T鎭_�|t�Ѿ�7�{j{�����sܡ�d2��	�N�,^R���/Wk�Z�Mzo�Gg+���k.��[.�E����,l�䆅;�{���m-`٬�Ӗ�\)�+��G>{��C����� �@��,��m/Z�7����������#_�~Wm���V�1�|��y������~��W5 =M�<CWn�r���ޏ����U
����N�,Y��V���8w�S��6��{o0l�䞤����-f�_y�Ж�4���7j�6@�^h>o{��7o��իW��'�O� ��E�\4<��}��o���9+
�N�y7Ɵ�ǇK#�s���s[??ًgx90�M�l���������3G�;�4�27�Ň�\��&{jwH-_;�s�;�a��k =K���잏�=_?:��r��9}٩CKG~���EË
'/~~��~��K��;����=~��U�UsV��ù�������-�w�v�?�S[ޫ�ڋ�~h�;���k� �$�p��x�o��Y������S��2���x���G����=��k��P�g罍�ǂ���Q�(6{y�;h-���W�3���{w�SOC����뿵��o��w��! �s:�X���WL�����T�dNYzJy*�K��?m�����d����k�k�ڻ��j��r��y����O�[�OXt|yNyv��۾Zk��1k!M;����KG7�n�x��� �)�g�tӺWV+�ׇ>�`hA��gU�C�z�r&d2�<k�S[>3�kgwyv�z�]Q���5V�YQ<n����\��g��ZV9�E�;�~a�W��Ӑ�&�k�\z����z�Ư z�@xk޿�����������p���OXt|)�`�\){��s�?}��'�4��F������=�|p��fw��q�+�)����K�r?ԋF���ze�H'�)��4�a�=����� ���`��ˎ��j��	�g��;f�|)s�ag-^|P�ϚS��;g��C_x苓�tn����{�������[˧B��E'�G�hE��+f/<���Z�W�-�Bknfn���M׼l�ŗO �'��D����l��V�5;������sV�=T�W�%���ZZxޢ畿��;&��n�o�
���B}圕���P������=�q���*�B%{O�|}7s�U��[7o��ݑ?��S~p����r���=����KO*wCc:�����x�m���������[�omn��<j�Q�_�=��b����H�s�]�4��H��8��7N=\ ��@�){?8vu}����G��(������9+gd�~7b�\~�P�Y��S�c�n�uϨo�}�m�j=�I�UsV҃0��P[5wU��+f���+�I'�c���W��z�W7���� �� ?f�ͣ����W����R��9w������s~6�͜����O����z��G�Fy6��z�+ۿZ}`��ӗ�V�����/<��o�c��n��5�	��H���n����w �$�~�[�8a�<yU��=�����y�sW�3\Η�=�����[q���~n�V�~�������S��/<�|��cK�L����[����/�}��&b#��픪���]���_�z��� �� SF7]3<Q���TB�8l�a����!�y�y�3��6���_�?���"�}���Y+Ϊ���l�� /<��<p�dw�@�X+�Z\��M=�� @tz�D���Uy��i(�1�-���r���9+�������ƚ�ɧ�m���Ǖ����{x�t.�^|�F��E&�QGz5W=cݭ����W_���t`����N�'�} 3�7�.=�r�#������O*�7&:;�w��Ώt��߳����ɝ��54T�ٳ�B%��#~n�3�v�ښ�;���׮ߴ���^|�? �!Ё�����~y�R�����\8{�YC�g-+�u'w�}ؙC�=p��X}�������=ɿm���ӗ�Q9l��(��D���y���|~b�9m�wB���4�j�=�wm�Í � Ё���}k�6g�ߞ�NϮ�=!��g�[u�Т�E���=��:o�S[n��~�53��i�_������j�����^ ����#.��qowO2���{6�^zU�h?O�A"Ё�5����i�=��/e.Xy�pw[���sV�=��?7���?����4�+��8w��m<��D��߶��Q���ǎ}h�O�:���x1p���e�Mj�׽>텇_8<�cwJ/ZX螕�{�ݵ Ob_m_w����+�^0��'_�tߌz�����y���w�L�뿷�W�۵�{�g �TO���\����t\��=������_0ܫC����ƛcIw�4���F�g�����N����*����{�������N��v����4W/W��t͋7^|�d ����@ټys������N�Y=l�0�}�?7\��������\�Ot�|��It�L���w��7�;�,9��Fru�31�<7���n�I'�/�V���Pz���� 8d:0P>���_7+ͣC�A�_8��>z\���sV�5tۣۖ�x͡����5�I�s��Ӈz���6�sV�5������ja�G?|����� ��@������j��[��=�G\82�=98������+�����&�S�<��������y+���z�ґ��ӗ�V���✽�	��B���z�[?��׾m{ `�	t` \t�EÍ��5�|�Z)_�\�����j�t��t�Yy����1i�;O�{�{.����z��s/M4':��u_#D�{��Xe���z���'Ё�0墫k�ڂУJ�R慇_8�k�ڟ��Ë�_|R��~��i��I>������p��+�\�w��'�������F�qr����.��� 3J�}o���p�4��У
�B��V���H���]pLic,�ne�4ƚ��g��ąG��H�Ezw�ݙ���lU'���&!B�����6_�?޹��� f�@�Zwj�m���ޫ[۳�\8oչCsʳ{�����rƲӆ&�������1��t#�S�^�H�es�V�7|ۖ�LT[��Hlg��Fho�z���#Ё�����*�V����v����-,���d3�!`��嶉Z�]���#��;&_p�=w&��������?3��b���.��k/��#�!Ё�5z�[N���[z�)�N�,���P��p9*\>=��It�B\���%���~�H�Mw�]��;�3*_���j�L�v2���[F7]��/�|2 0�:з����������_:jޑ�0�����<��ʗ�}���������C_��n���=��ˋ�,8&����E7ٽ�i�/�v�c�� �N�}i�-�]6��86���+��脲$�A��/:>���{��ӽ��·爵uؙC�y��<�I�}��ɮ��v�L�X{���������� L+���+n�b�����4�2/w��3z..��	��W�����m&��3m��P�R��O\|b%��L�d�^q�Ч���x�U����NH����_m޼��W�6�`	t���˭�w��r�1�|��Q��΁�Yq��Ӈ�ݳ�~�{w}�1Rɮ������t��9�����D�F�衕k-�����S�	 L���5�_s~=_� ��\�{��������E�͋��b�]��\��];�V�������=�Z�{kA��J���b��Vn�����o�x�c�i�3�h�d8�ew;f�1�/?�2(w�?[�B���?�����1]"�I���m_���#_<����N4&:������X�={���/i�Q�����P�X�˩�� L���X����1�������9+�:�gj^e^��e�}e�W�����4����/:�#�C4�=iZmLv�N�������2�w�W���������q�\sg ��@_X�y]��o��5@*���́�}3c�T��x%��Wۗ|�o�NYr��t�\�N;o�'�~�c?|�]��i��:��1��? :��N��v�=/��r��9w��C��́g��%�/OL��#��������[�����+�8h;U����7�'�kcI����}I�5�	���=���_}�k��5 pP	t�獾g���r�7B���p�ag�r�������Y+����OOL��@D��]�]�_��*=�Yi�]�O}��v���K����}Xa��ݰy�ǮZ}U3 p�t��5g%oOB���S:~�����Z!�Ϟ���������a�[��N�闷���#_0�T�V���tj�ǚWL=�� �A#Ё�v�M�g6��sC�
��	���7b5R�-Y��՝���'�g�wS�����t�W꯾r��z��� �@z�p��{�Z�b��9{ř�aUΝ?Gͤѹg׽�G'��{w�SߺoksP΋O�vH���[��9 pPt�g��u���)������J9_�7b�I;�=[�켧��m=�I�4��^n�����5o���� <g�Y�|��ǧ���UsV��^��gi�?t���m�o<��z�]X�$ө����*�e��L�=i��ֿd�P?�Wf�U
��)�Nq�������}��w�ƚ�Cd�����n}�Ƌ7> xN:Г�#ɕi�����"�Y��Y�N<#�N���G�U��M��!N��)%��?O=\ xN:�s��t�/W�c{�׎Zpdq��BW�=C�M>ֺ��j�V�vv�\�T���7�u���yێ ��&Ё��n���yw ܉�N�X#it���7j��ok�'$�S
�ڟM=|c �Y�@OY�����G�q���*�l�'�L��T�7��qw�tv�=�R�������x�;� ����V��3�3��,,Yjk��^���ǾS�����I��Z��;�}m �Y�@��y���������K�ok���%_���ɱƘ���㪅�/_r�%�߽��c�gL�=#�t��ʽ�'-9�\̕Lm��[ڻ���4���@'����d��� Ϙ@z��{F��U�	=`nen��yGO)�$�;���Yn�j���W�^�:	 <#�	�Y��NH���.�����yR�)�_����=�=^�Cje��P��k�� xF���=��,6)���*.Z��)��o~��z��9��F��� ��1/"�����C5��k�L.s���O��GZ_�����������lZ�+���� 8`�چtCv�'��F��/<�T�W�{��}��_��A�à�T�?��N�<���&/n��ȕ���1�.~B&���~�����o`�4�׿o����k�	 �D�Ul�v�'->������I�]�]���P'�ٴ�y��õ�"Ёh]v�eG�&���]��[5wU!��������0����Kn�����_�zW* �D�]��Iw&D�E't�Y=��4��W���@hg�Y��|o��� ~&�Di��͹�
��B�����ܲYK�F��@7ο��+��c��9�V��=�$��@�tG���*���u�UK��?!��C_���!΁i�'u�,����~ �i	t J�r�������Ë�=?��~��w��9�ӺG�Z��uS� <-�Dg��F���UO
�{���\��C�������O�Yh�tC��-We�� ��@�Ӟ�yC����V��/v�|ʃ�lܳ��F x
�\2w��c�q��� OI��i[�"w��畜=����]��g)��:���@Tֿo�KƳ��!b�K���f--������������A�7�F�q�%7\2��k�= xR�JRIW��������^o�;_����N���	i!������} �I	t *�|���R��Y9g�@On��F�n�xFڥ��)	t ����_ޟ�77D��yG�2��@��}�7j�����j�'�yߚ�7��� ��@��ʶ~+D,�͇#�^l��m�-{��NxV���gr�ߝz�_ ��@��!ݐ}�㻣�޾r��b1W�����4VK�|�.ہ�$��J� OJ�Q�����s۳CĎ�����'�v��m_�L�Ĺs�9i�'n�䆅W���]�� Ё(�C�+C��V�����s�7�Vm�9�	 �Q����D�N�w ~����������'v�"vԼ�v�|Wug���8w4�b���.�~�@���>����H�3�̊��2�۝v���w��`g;p�r��F7]3����' ?"ЁC.
/[5wU!����j_{���Z�fk;pPu����/�zxk �G:pȵs�����r W���u��V ��B��A���R��FO�+B�F����+�r��������wW�4iۧ ~�@���e'���-�j���T�����켧�h��}	`�2�W�r��W_t�7 ���!��/[9gE!���D�e��� 0͚��+��� ?$ЁC�׫�>)DjAea~�8���G�^�I �n�Br~ �G:p��zϾ&��^��b�a�z�����c����h��]t�E÷\~��� �@�¬ܯ6C�2Sߖ�Z:P��I;�7�f= ̐NH�.�^��� �@�V�}f������r����p���7��Iw�3���� �'ЁCb���G�
�:l����{����|�`8`�%�4�Y$ 3M���xc��B��峗�������h��Uf\#�\�:��P I.����9�J�20�����!��Nnɲ�/�z�?����!�)$��H-Y:Pύ߳zbI��� �:ph�r��C���,�v���f��A'�� �����-'�e�Fy�y![�t'�����9�f�q�tC���Un� �@f^���!RKf-�gB&@��{{�X=�$ө�_����w�&Ё�Φg�H-^<0ϋ��h�[5��@���{�@�����.���Z4�p`��칿 "�ʶ� n`^�q��u�ζ�����Pqh ΟO6&���]� �$� �@f��ϝ�l��ґ%�e���4��ģ�K���7�����1��50/F�H�g�H-Z0ωݫ���`+ D$�ܖ�[��F� �@����C�-�����n��"= D&��wϡt``	t`F%���!B�|)3\�B�n����s Ji�sb `�Q�\�<Dh~e~~*�����f����ɠ8`�	t`�\z㕫ja�P�Ђ����޾}lG+Ma� Ћ��N�o���̘����Z�Ӽ�y���o���V����4�x�� H�3��&��e���)���@���]�v2i&=o��'� ����d�cB�*��l!���n����v�t��f�@�@fL'�Y"4�<��Wϻ{��v z�LzD P�1��Z"4o ��w�N�����v ~��$ (�̈u��U&Bm8DhNyv�����v���@��l{a P��f��P���٥�}�|��nu�$�� J�3��vN�fra�8������N��$tJ�Z�@fD'�)u��G���$�v���/	 =�����������ȥ+B�f��{{w8\'��@��:�N}w[ 0�I6]"4R��@�5���v��t�� 0�:0#�\�(DhV��}om��s����a` 	t`F��N�Sy+�J���Ƙ@zJ'$K� ���ۼys�_��
i��P��'��۵N�݈��<�SK��� 0�:0�>߸{qZH������V.��:���VρޓC` 	t`��ZQ�+ʙ�Է�����t��tBR	 H��/Ӊ2Ї���|��s�%�SZ�y]����� ����2QNp/��}���VЁޔ�z�z�-`�t`�����r����ۧ���N �A�y��$w��L�N��*�}��v=�Ёޔ43�Z�@�_.�"T��z�{�ݰz��l.�  �L�N'�@/�J}��^k����4Ӊr~	�t���K�aV�P1��g�k�t�g����(��$Ё闦��B��߁ު	t�we��Ё�#Ёi�	i!D(���{�����L1 �L�L�*�|�ࠩ�������O� OB��.M3Q>���
z�Ӷ���N6�����E3�g�i��5�l����@�f�8Q�h�M�[�s�l��%椓��?��2^���0����=3�-�~�ǒT����A�@�]'Ms��p&��.I��g �̀N�+衯Wϻ��c�Yi&�u*0p<�Ӯ��l���|*��zWR�S����vS-��m)7���=������ui?Q<	�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �  O��h��2��s�dB'_�7 }O� <�N'�U�M.:��C����Z8�� @��  O�X)T�vy_c�>7 �4�  O�2����$�V�5+ �4�  ?�М���B�J� ��@ �2�����9�k|I'� L� p 2�Lgd�T��_��i. �A&� P6�m�~lb���p��_��t�>��!Ӫ�*�\��ods�d�~�����]���5 ��@�S�f�8�ora��� },_*Lv�C�ɟ��k L�Ї�Fyb�Ĝ`.}._��F��:?��� 8�:@I�N�^�5�-��{�B�><d��\���$��D�jjSq` L�y�{�Y���C�y�~��I���� �F�Vi�g��\�5<o*γ�N���� 8X:@K��|��������L&��̟��LMl?P�_�`� =�QkTZ��-��n�/y4��F�O认O}��� <[�{w%�]������^�{k�eyw�Ƅ�!�d�K�$d杼�eN�!!���cb�:���[��p��c��wf�aBl�}1�ٖ�Œ,����.�����[����ߪ�]tI��������F�@]�ͨy� �BIdF���닅t���\uq X ��jg��Ec���xq�K{m���s�I�5�@  ��@�0���Z#F�s6�0^8�e��X�l�hF��� �t �ǧa��F�l�!2q^��N�~�  V � ���4��H�D&����j�թ�� �B���8>�.[��g
��X�6_�Z3[  +�@ �p|�]��l)[K5ʍq�� �F��%8>I�R���܂X�Qi��� �t � ǧ�EIƫ�
sb�f�Yj�Z� @�� �G����fa�8+�j7څ�bsB  �" ������l���y�8Y�QJ�X��������  �e: �ǧ?�zn�8Q�6��V��/Ԉs @O� �C���r�_0q�H,��Lm��J��
 � z��ӀQJ���Ҍ�P,��tu�8 �� ]��i�s(�
��c��b�0��\m�h��, ��t �"�O�#���D�r}�PDn�Du�֚�  =G�@�4�<�?FƋǽ���H;չ���g��  }� t��� K�8/Oe��X��f�<Լ� �  t]n$7�ʦb!s�au�:!�8 ��@  ]�-f�3�LU,d�f���+ �w:  �L1��-e+b��|u*h9 �:  �T.��+e�b��B}2hy �:  Xq�l�Z+̉���x��.
  !� ���2^�0^8!�j,6G[�ֈ  `  �7�6��Y�T��,���1 �B:  Xq������D��ڍv��؜  ,E� �eS��Ek��o���B}J  ��  �E9*(M��?Gb!�dk�i �r:  �`J��8Y<�*� S���8W ��t  pa�D��빁X(��Tu��J�8 @�  �B��xq�K{m�P�^�Du5q H  �/]/�2^K,�ڭ�q��v �!� �yɏfS�TC,�#�,����?s� H^�  �9ˍ�N�s��X�糋�u�S @�  ��d���L!Si-�:W���(-  $�  �*�r�����L���8�0+  $�  ^P:�^̍��R���d�r @��  ���L���ω�j���� �@� ����^�0^8!�jTc~�/	  �@  ���Va�x\)�b��bs�Uk�
  �@  ?�q�vq�8ck�7��R��  �  ��\�'K3�Q�X�Uk���	 ` �  �C)��s�U�X�o��F�1)  (  �u.Qa�x���@,䷂lm�6-�g
 ��"� vq�'�Ǽ�닅�v���W�s ��#� n�8^���^[,�W���-�  0�t  ��.��{�%
�ȭ�V�h�] `�  ��H�D*�j���P�չ���9 `��  �l);�)djb!i�6W]�C�  �� �����bvQ,���j�a� �!C� 0D2�L%Wʖ�B&�ks���3 �"� �l���͋�j�թ�� �!E� 0��W/�N��j�ɠ� �!F� 0�ܔ�,�g�R�rc�o�E `��  �8�[��ҌR��B�Jc�Uo�   � T�봋Ek�Ym�Z�֨  � ��tF����0/4�  �E� 0`�Raq�x�qU(j7�|�Ҙ  �ct  ���ǹ빁X�o��B�8 �4t  �N�'� �Q�J)qG�R��}�׵�A+��檫ļ�   ��@ `0hIɂ��_�M�+�v׉\��&�ͷ�c�w'�v����  � ��R�,�j���E��9<Ɂ8�{�8��}^����x�Ы��V�~��  ?B� �t�T�8o��C������n'��h�繑	y7�|�ǋB�VOTWk�]  /�@  ����S�^}�8ޝ�ֹ�;K�nb=����#�,����?s� �9� �����y],�l����H����Z�xge<  8':  I�J=���Hk��q ��!� HG�*�,����G�8O  8/:  I�HK���XJ��Q�$#  ��  $��v�b�8�G�8�
  � :  I��Wieo��Q)��  �F� `;%��q�u�r� ��  ,� ��B��\QN)
  X6  Kiё�qM�Gb�Pg�8  �"t  ,�cf�\��b�Pg�v4��  �2t  ,�l�;*�0J�&� Xa:  vѝ��勍"���|LQ�  �8  �������b�H{Q;"� �  [xb�)6���q>�D9  ��@ ��S�⩆XH�8Q�8 ��t  �͕Z�u�Q�����b~�  ��t  �ɑ�J9U���J�zL4�  �/�  �#M�v*b)�[{�)  =A� �J�q���R��8O  � �Ӣ}'�,���8�H2  z�@ ���q�ϋRZl��8γ  z�@ �wB'��k3�n!�GE	%'  �/t  z@��ܬ;�y$6
t!��  ��!� �2�N��8�A��@�  ��@ ��t�Lk%��(��8�G  �� @��8Wi� �
�F��D�hT)%  ��t  ��1眻�-�a�_�s  ,B� �*�L���F�N�S�9  V!� Xi�,�q�Eڋ�q ��t  V��TU<Uiq�8W�  �!� X)���8�������s  lF� ����R�b#�U���b�B   �"��K�`h8Ҋ�"6��\�8׼� `;^���0T:�؄k(i��� �2���q�$VFN��빑  � +Ik	�� X�;��*�,����yZ�h:~^�.���L:�峁  � +Č�~�D�9J�8��E)+W3�q>*�d��j{a��|�g4 � + ���g�|��Nƙ׶n5��8γ����2��l&��2����!�`9��v�w#�z�a�EGN�5qn��������V��u�B�wŞ� 0 t �@Li>:fF�E�	l�8��Ϭ 
A8��j�Ly�R��o �� �)����8w��ӊu��8/
�JiU�֙� �@��`vS���>�tg�vG�b�Pg%���2S�͌�|1ϔw H0 �Sڇ�J����-6
uF�zT0��0�Ly���� 	E��9�@�A�
��'�8�[b�H��v4���$3�����g�t&m�^	 �3#��,̨y�z���ʢ��(�^Ԋ�u��hԛ)s$[�K�!��L8Bm�)OU�Su��7j�xa�V�s�� 9t 8֛7e��S5�P��錜�bV���u��B�u" ,G��s�8o�>�͇�#�8��B�8oFb&��s[�Dz����r: �"���'·�#-�v�b#�U��cB��h��y�I�<�ڬ�x�m���Ͻ�o : <������v�b�8ε�s-)��lgFԳ�����E:rˡ��{nx�3rϧ � � 2q��
���1U���b��-�_;�"Z9��С�ƿ�Q|k
�IV��lyZkI��:%����[���}�>�G�n�S��:mqTg}�2�ۥ+79��{�7;�{r�%.��û���+�|�\�����'��ͷ߲��v~� � #�/�1j �W��/ҪPʷ�r�l;�T��ݷ��靯�i��? \(�P�Q��s �.�Z���#�#����>�G��^* 0�t Cǌ���q '�JOJ��fg/��w�������� �`�t�ZOy�&zC8 XI��t��w�W~�����O���g �`h,Ź��\���S-E�Y�������Փ�}�z�������� � !���q^K�!���LL���֏���}�q�k���I6�0Ht Ϝ�{r�8��Y�t�ww���G���o�w� :��W�6��S  ����ި5R���~<3��n���y�=$ 0 t �\`�M �s�(�s���SȵҲO?uۍ��ow�s�n��#�,�L �i�ڞ�0.��X�a:t���#�;* �p:���l�<� ���ly��t:��R�\�������>��s� @�� N��v��  VD��L9�������e���o�o|z��F  ���0P� t̅�  V�9�0Rl����BZ�z�?t��_��?s���"���Y�:q ]W�j���k��Y�n�V��y�K�3���"�3�c"]  ]��2GW�|F�L��տw���O���_ $�` ��9� ��]i6�ugw��k����]����ol	 $� �ر z������v��Ǿ���� 	B�H��vl��3r��ٺi܌7{�o{�/|�}��� @BpQ ��z�F���p �'fyQq�`�zt�z�q��6. �:��2�l
 �c��0�ŹB��r���z��?�W�_ H @"��-�lT$ ��2{�x)/J�SV�GZ���p��o���?- `9@�Ahvfj; X��hzf=��8N,�Cw�q����� �#�$��Z�:q 1ˍ�պ���Od�.���7������E �� �Yo�� ,d֣�z>�vD�陿��N	 X�@�fj;���̱�f-��G�-f�o��[?�{>$ `)@b0� �g��kJ��������Z:�D0�&�� �3S�ۭ��Τ��ս�mg^��������s�% `!����v3mR  �Ь7=/��rW���c�v��o�����i�Zy �����  #�re��Jy릺�Y?����U|��	 X��^ V3�$�tI $JN����"�̌���ۿ|�o1��6: k�5�Lm��j���h�%�ig|o�?�O��_ �� �ǹ��p �\�9���ʱ+ `���02u<G@�ٺa�E��?|�g��>� Kp��J�g�� 0ƙQ�|ֺ��ǂ��W��@`�u̦Bfs! 3#�Lsw]ǪQ�F��{�mox�g��� X�@`�f��� `дM/_��b������O: +p�*f��c� `��~��A��kձk����������/
 ���*����2;�缜U����)<��] �ϸ`F�`��۾��f�֢�y�o����w�Q �#�5=���n��\!g�Z�������_�w] ���`F�`8�Q�L.�v.��,�� @�� ��j�y>�!avt�m��k�x������ ��b }����s 6��k%2���� ��@�wfW_ ����t&�E�vr�W:���/�t 2�f˳-ЃL���m�s�g��ُ
 ������y��� �ab����^ʳ�\�rP}K��@�:��j�=�a�}׶@��� }B��09Z �������}�{��������� @�� ����  ~��d��֢�Go�?� z�@�7� �ہk[�W��Z�> ������  f�SF�uk�������7��?��� �!@_���  9����2��B����;�{:��"���� K̬*�e�&e�x� @�� z��� �S�i��u����^���?}�����y�!����3z �q���=Q����}� @�� z.�Y �q6��^���	 �����N�Lo <��段��y��Im� @� z*ds8 ��A�x)/K4�Vn׮]�o��% �:��
X 8���@מV�?�÷�w� �@O�)� �i�x�Z#���� z�@�3f�"�� gb�qkuin �@��^�9 �E�k��x�zS%�!���� gc�:� �n����w�Q �2@ϰ� p6f9�XD�?�J����& �e:��0g۲� p6Qd�r�z��%!�� ��'�0�jD `'�f�mo��u�2� ��� �Ud�kF��q� ��DFV]l �eۛ�-��
 � ��'l�� `/�,J�=�z!�� z�' =�5#� �scf]y�+��<���'o��c���# ]D�艈� ��䛺��Qo�_"�t��뢈�s ��뼩kW�K$�K ��@�u�� �W��z�hF�u ]F��:�: �<���ю�	�.#�t#� ���D ��@�u�e�� �gۛ��9�.#�t�� Ηm#�
� ]F�  �:ZGb�8�S ]F��>-�� Ώe�Zi^� t���"˦) p��� ��@  �ul[��:�^ �t�f�8 @�� z�@   �®�| ��@�.q'�t���*���s�����$�!d�wa@� za(/j���������J;AWān��P���5@��(�Ȳ�2 `;M>:��ӌ;  �� ����:#�*  Αm'�(e�O��"�t���6 ���w C�@�}\d ���7w`�� �����U �|Xw� � ���P;�  p�th�1k�A�:�����uy� ��0�
t ���t]E� �KV:#� z�@�u�� �܅aH::���) �Or:��C��:� ·#�Q%�� t]0M p�t��ۻ�t �@��	D)�9�  p���2:�^ ��DFi�@ ����F0�x��A���O9 ��k��V�`0z�W�z�0��8г�  �&���@�+:���}��� g����5 Ê@����#툣" �B?L�et �B���Q��M �� �sw- �u:��	�~�M� �3k7�\�Z<���+�)d �3i5[V]�2�@/Y�`��]nIk_�0Q �<�f���%�@�K:��1]Q����  ���jg�2��!$ z�@�S~��dt �i�-��� �Gt =�j�ҬC ��Y
%!�����ڭ�#�C <����m��L:��28�fݴ�  ��n���^u��sF������f��.� �g5ꍴX�(�k:��k���h�i� ��(ӁXU��9�~ ���� �j7�9���t }�4w ���s�9�~ ��Eg��XQ  �-�릷���@_t������`��M?��9f@/� ��Yk�� í^�'bz;#� z�@�7�E�W+��$ ��	Z~.B�ʗ�� ��@�W�z��)d+ :�j#/�a�@?� ���X�ā. ����k6��X��s �D��+3���� `��ꭂX�@�O:��3S�% �H�Z�ns8���7@�5��8VL��| <���0���]��3�9f@/� �P�Ԋ���  ^�R���s�t �F��B�ZO�KyO�N  ��4�����[�}���JC� ��@`�V�U̎� 0����uG�/4��`t@/� �Q]�����+JB ����l=?���:��#�X�l�Ӭ6�q�� 0pj���G��m�܈�)� ��@`�j��ɕrN|	 ``�~�m��֍��2��D�K ��@`3�ި4FX� ����X�ms�%��:��#�Xg������� {n����Lo7q�@�� �T]����9 $��jq�b����:zn�$ś� ��@`�F���J���r� H�f�Y
���-��u��pD� ��@`���Jql�8� 	��ȭ��Y�����)IU ��@`-sV�Y��ʦj H�z�>b6������w~�x,��u: �U�����S�]�d��0S��Sb��=7�*uT ��t V��HU�����  �2_)��.$�S��G ��t �3#0�B��  !��ƈY�$2q����Y��2� t� *s���ꉖ�s1# �CQ�֍��]{n�����X�G�.#�$B��Qi�fGr �Ve�2j��p2��H�T�s�κ @�� c�����3�9�E j�Z�v�m��v�BFύT�j � � Q�s呱�YQ��� Rfj{e��K]h���5 =A�H���b��� `����M�.tz��v2 z�@�8f�{*�ʻ��� `�f�16�SۗdU�� =@�H���ɵS-Q
 �o���3o��������v����� �$RER�]5�� }���-ϕ�b�厞{��z�G�. �:��2�)[��h��- ���ձ(��7<�E&Η;z^Ѕ� @�� ��Pɼz���Gf�ں9 "�i��\��t-wc�%y7wX �Gt ��zt�l�RH������! ��[A޼A*[���%Y�g�8 =C�H�+6\.f�|C~}�:U��>� @ט���g�^wnFΗ;��0�P*�?* �#:��ɍ�����a�K'.���-ΰ�; tC���c6/)2a�b��A����}� =B�H���_*���a�\���}e~�]� ��*s������X�87J�xD ��t ���2rњ���~�wݖW�ܷ��r�o�;� 	�(��Z���w]뢕�ھ$�
�
 �� �.^w�xn�Wan�d~j�u�/?q_5�" ��]k���մXl%��w/~�-��/ �C:��q�#������y:L�_��:�/{�G:K��B�M�P�/��r+�F6ʶ>��� �!@�l[�U���a4���|�����8���|�~�]��/��L����vcT� �1@�\���s�qZk5��,�d���w>� �9��03?37"�3���m����?	 �� Q֎�����9�DQ��f׌đ��{�{- ��9�|nfn���Ԍ�^w���JOMn}� @�� ����c�Hߐ_?��?<�`[  g�ŝ���=΍nĹ1���|�-� =F�H�����_wA����Җ�pmP~��n" NC���0�0��g��Xw�d��{�> �$��.��\����\4�}Tk)?y�I_  ?��5q���qޭu����Q�V�> �$B6���-�q�H�E��G�� �0#����1rޭu�KF���;�{�a�> �$�9��u��p�H�6�m4~���+,���4����^�����( �': 빎+��xE�Dzm��ϗ
u�!evk7��'������� ��@`��I.�[�� ���B1��L0\"��8�֦pKF���Go��A�>!�XM�����k�Ƒ^]���BS	 ����3s#I8J����Wc�U ��t V+dRʍt�kDQ���8�[�uB������|1)q���O��R��׽�͟�O
 ���j�fU��}�\��:�@���I|���q��Hw<7 @�Z�T�/�$!��c��&dr�o��o7 ��@�uf�#��=���A���r��?���b�Ƿj��)
�M���`��j͑�|%+	a�ۛ�=������6�>#�t���"-˙Ny`��8ҿ"?}�Ou5ҍZ����r�ˤ� I����kc�j=%	��87F����� �3@O�� ������q�K^��H�7�t8�|���U� pZ��ly��jw�
�e�S�� � ��gV"ҟ<�Wځߙ��:nW#����0�R�c� $������HR�Q[��8�D�`�+��@ �:��2��M�/���އ�W_~�v]������Rͱ�;�$�~�|b����ڗ���皒�w�f'��������.7���|��g����^͙��1l�\�g]: ۵����B%#	ӏ8w��G��o X�@�s+�G��?<G����T��Wuf]z&
�l.˺t ���S��L���D�77��ƴL?�띻v X�@�+�3�����������.d]��k��n`֥�Mqԅ� +(��l��B)i�͍~Ź+��p�~S �":��Y�H_�����E�٫~FO'�~���Z�,�
�B��t }����Oկ87���}w��� X�@�W+��v]������5z�誮_�)��Z-�Τ�S���r�<��)�F?��%���
 X�@�w�-�J-��VВ/����\o_��'W}�V�� �/���@τ� 7|���]ڗ�3΍�h�Ю��W �2: k��9�a�W���ke}�֫�W��(��b5����T&�N��2�D�Z5����Ŵ$T��܌��έ�} � �����>$�ͪ��%���Y�'���]�SA����f|�I�XQ�f�s������������#w���/ X��ϒ �+������ުɫ/�^�2��\����e?�h:�cFͫ͑��b��6_bK�;��jw���X��ϔ p�B.C���d6S9.�み�W_q����I�?;���n.�kq���(�pb!���-qn��5�����Y �Rv<[�i������H7;���ү�r��rӕ=�����	*�9F���57�y����R��M��y �� �f.���M_3]�������~Ŏ�K/֥w��0���� ʖ��%��'v��0��&�m�A�}��oz� �� �g.�L�/��t��c{e�� �_~�.�J=M�+��L6f�i�M�<:��z�>R��S�p��y.̶�\��� �� ��0����nw�:'����C^y�+��U[z:B�j6]�����y�M�� @̯�K��r.�皟��Ǩ��w��;_�s���@�� c)�Wb�w?����ˑ�#�'/�Iq�gW��֪V��S����e��1stZe�b���3�|�l��T����'��w $�}Ϣ p���)ơ�w�:_�Ǐ�錨�����#����t�d��\6�ҙt+��f Ι�^���k���nشܩ�H�Պc� $� ��
�r�ů���90�Բ���Δ�k�]�/[iO#�Dy���Z͖k��{)�'�q����NV��R�C���0���]oe:�a�z�S��u_���w�� @B� +���\��ç��=��i�Aȷ����;����:ɥs=��i�㤲���q��'��0t��f������r>B�h/���͗�Bc�u�V  At �_�m�J�J���G�����sOwFӯ��z����_u�Q�����X6%�O.����|�8�̗�(_:�FN��1���l it a��:�K��������x�����n�?>�O�ez�~Ŏ�I:����Y���\:���L�L` ���(]]�����}�������Z�W�`�;v}V  at ��-��^����C�ٳ���|�̔g��;^�7Nm��0Q��v�[>�N��\�͈:� �N�ʵR�V��,���/�E���э� H��{� 0�<�U���:�0�^�K+h-�������_�k.��n����]�������#��p��>�}��k���p�η�\� �'� ��U[��ȴ���rt�زo��'���ayɶk�����v���L:�0������y�Qo�uU��/Y-���;>�A��� 0�قz�^?rh�|���H��7�l֦�ѯ�����.����}�V��Ʒ|'�3��8�u��T����:�>����=8q�� J�%Ũ�xю�� H0�@3��_��rY5����{�QY�c:qH���+7^���t�]�w��ҩT��f��uB�5��ʺº�ֱ-�B��ٕ��/�9��}ߗ>$��D���p������Ϳz�`�S`h$� �azdJ����N����#�w/��̹��?�90���l�O�գ��:���}'�e]���l�W�j��q�j����҆l�����w�uͶkd�0������>��Lg7�ړd���_��_ H8���\O���ɚ�5�����r������%ٲj��v۵�����av�Qw�J�r��Ӈj���f�:p!�sc���5�5)�q_�������DqB��{Wd�N�%m�|�T8u�����. 0 ��, ˴ez�Z7�V�o˞#O���ū����엃��:�ޯ�t���B��"��Xz,=���b��H�H}ω'��V�R���ܦҦ�xn��v���
c�����ǿ�9�1)�8jnd���J&R `@� ��9.�.�N.Z�]�ѯ��h�Ҵ�'g��5[��[�6K�wW2#�*T޺ܺ��֗��f�`�Pt�r\/���)]�T�QXi$;�n,�/�-�M����j�K��/{��,M���g�$u��p��[��o��w �|F��flMgm����C�ȅ�bcQ̆t�����/����%Q��dnR��n{u[�^<"�O�v����*r�n6�l�VZ�[_Xޣ�/(.�+7^a����?�/+��f�%u�|�fgӗv�s�= �@0�����^t�l�ޤ���We�^^�ǝ]��O7�����H)W�$ԣ��ߓM���et��ԏˑ�Q�Y�֪cX�.N{K�
�Ң�k�jޠ��k���w��2S�$�\�3��|꽟|� ��!���GW�׽�u����<ԙ��\f��������t�m~Q�7�;Ui��N�tnZd����q9\~ZNTOH?���T���+��o(��潼��ރ?���������3u>ܷ�[f:�	�k~&ŰX[�Yu� � "���㪫��X.^��s$ۓ�����F:�Ǐ쑽���%�.�Wm�R2��5Wɝ��������X��Z8,��E��s<���&���67���L����u"/�6Q��_}�k=?�mF͍t�
6��^w���	   N��)��/�i���7�ƊM{7��z8������ŷ�͆ub��)���e��&�9Z=*��I���n�_�I�u#k3k
�s��c�Ė�-j<?����}R^��2(an���[���|�-w�P `@� �֍�U���_֏~T��=�CE�<��PvǏ{�K:��Ie�6AJZ�eSi�l�"�vE��sr�rL*����UH�Ԛ��tn:;��H�Jm����1���~���׵��e:���b�����c! 0�t 8�q�/�-�6�o�����mlvP��S�#�w��kv�s��zU�QER�R)�ֱ-��~'֏׎˱�L��CzE�S�)g*7���MeF�#^���5E��w|�<��C]����~:���o�ݟ�]�G��92����W�L��Γߑ��V��zT�f���kw�e.�b�(�2���f����j�j���b�Y?Z>*��%�JK�)Y5�J�S2���ԙ^:y ��?�Y��ȡ�];rm����j2�<������ � � �i�ȴ��*����z��2_�_��6k�M��~�Q�:�E��p��TJlfb]���c2�.��Tʭ��Ʊ>W����\g�<�B��%YU���8��sc�<���J�I-��w��=�X�޸2ann�2��T�z�|펫�^�F `� �nT��/Hy\���u�߼�u���O�w�>���bfTp�̾�m��*�j㕲ab����2����ݼl�$[ƶ�ٟ��We�Y�c�ǜc�	��3Ȧ�2Y����L�$�������+����̊Y�#Og�֙?W1,�/��v�Ϳz3�S:��[�[�#���^� &�0V;�^$[Wm��-�u��|%͔g���,�q�t�%�}ն��<O��3��Y��5��l(��+O��Ͳ�9�:V9��ͅ!#�C��)�D~\�� ��OH��J�(�m���c�և�wf��?ڵ��=̍�ε7�ֿd�n� "ɸ��hw�|�ܭ�n����'���� ��ԋ6_%�ۡx�Ay��c+>jf����o�{�'�M�K�^,�\I���
/�xyU��Bnsa�V�D�Vşo-�q��N�f�Z���*ù2���f'
2��yJ�N.�xƩq�A�wfҘS���a�|i:� �D�p}{���ڹ�1�!C�����C���;�{���7[nk`�{r��z�E/�m�	m6�z���+v4������q>�l�� ���D֍��~���DQ�$�h>�����Ƣ��Ӂ�r��[��\m.�k̇u�=q
�����d$;"#��7�O�?%y��\uN�)�{��]���07<�Ee/��;�sǽ Ch`/��烷|�{�?xݞ`�o���m5|�l*����b�|�e�P$�镞�n֩?5{�s+e��c��h�E�K�$��1Ym�7�48%��*�J�M�M�s]�k?4#��v�5W_ˍ��֪�$l6��ȸ9u`$7"�TA��b'�Sf��)��:J��-��@gm����~�a
s�ю��l��Λ��� C�@�Sw�z����7���O�m��:ҍgC}����Ïv%ԍ�fU��=���tF��Qm���%rT���({ی����#�H*�����f���_�G�v=�������F%Zl��Jk1b#��ȧ�R�$�	���)J)S�D��1n<��IfF��yB�������S[�n�;����[�[ `�� z����}ۇn��=����?�nd��N�_��2m���>�hW�\2Ǚ�}�s�g�}����MF�2HL�G�D{Z�^����
��;��N�
�aկ��v-��5��X��vM�A��(H�@nW�ݴ�ɥr��rq���x!��8��q�ɑ���%m�z��~y�ؓ&л���1�3r�=����o��� C�@�w����f"��8��C�F�3�~���������>��Z�����zgWys���m��vn�TFճ���)�+�bg�W2f�=΀��C	�fЊ�a��A+lFM�L���o�,�<�#��J�MI�Ku>g܌d���AnvO7A��o�r;���Kn�~\���0
����c{�����R�n�]�����E���|���?   @��H��7�֞`�_N0TCF��v�g�(��=��������}=�V�ܾ������[Wm�L���H�x7w°3�'�Y#�.�O����`��V��a��~d>���{a|O���#hK�ݔV�6?.���n��rt>�s$/����S�
�vMx���_^����H��7��'N�:o3~���	߸�Bhis��ޙ}b֗w{
�����as��n�#��]o��i� �@_�z�G?�oj�	��ۖ����%�|����������&�5jF���As3�!�t��'�wFW��٠.��7G~=[Kf:w�|�����9��DU|���7:#��~?���8�M�ǱG{�=~�����i/�Q���2��3��)���ک�~���?м�b��I9)e~�\'�>�R�g���I�W���LD�p��Y��}q�?5����޳�m�܌�3����-�� �Y:��3k�o��������o����}��Ҥ\�O�K�]#�-Oy�+�ԗ�s���߹��3#ꛦ6ű�n�F�/�	b�K�O��?�3�'�.vX�磟Q>���OǍ�h���mw��n� ��@`�]��u�w����{�o�ʹ1s\�9K݄�����ӏuu��a�p6#��fFi׎���q���� �Y��3Ǣ�?��̑C���=��ü��tҒ
���ް��]� ��� ��?��?p����߭���9���L?77���9����꨺aF֗����X=�J�Ol��e�0&����>8w��G�87�{�i�ϗ�2���E�t׭��  N�@`�]�ܵ��߾�棏��
5������t�K��/�٨�a�q]8ֹ}w�w;��f�����ck� �e�g�������Oˡ��2�8חc�-?���7�8�^q���  Έ++ ֹ��;gv�ڵ�[���9�f7�u������އ���1PK�ͪ<��c�����ℬ[ۙ�zt5�k�3�Ƣ<�p�3}݄y�v^?F�_�x46�Z�/���w �"�X��o4�7��}o�����/����+��y�@7GfE=�0�|]��=x�α^k��tF��ı>�tx��F�.G�f6�����f��?�a?"�\M�_���mozӛ| ���j���3/}����~.�Ô�$X�Vkn��uì�?p�@�fdSY���U�6�J�JS��㜙 ?V����L帔k�L[?;��;��k����}�e���[  �@`�O�㓯}��r׾h�[C1\���a�t
���n�K��i/݉�8���ȔL������F��W����	��c܌���@�Q~��_-�,�ۧ���+ ��B�H�?{���v�o����M���s`��L�7�F���Y#l6�2���/�ɏtb}�4�9���:.�>��?��zYfM�wn�2�y��9����Yz��ǋ�h���?��]�Q  �@��޾�����_����ߍ�Y��SG m�u�LW6�fnO}��}�rd4?�'K2Q���ℌ�%奈�2#���N����;���|_7t;��(g]���G�֖Ԧ_��ֻ8F .� Qv�e�7��u�ʣ����JS\I�'c}�E]
9���nF�ق6��渹��O�w]�����m�Q�J�r2�kq��!^��m˟��a��ʙԓG��̕w��9 \0@����;j�o��������^��r"��'��`�vs���:q���7�^��}$?"�숌ƟGr��6b�>�/�?+����#�^�J��	r3��X�j��a����J�zw�7?s�=� ��� �����/��#7��[�o����v=FS���-��#�&��Q['��z�����q�u�R������/şs�Ph�g���7Bj�ڳo�,>����0y'e1u�{<�F��mw~�ֻ�. �A�H��n�����p��,��W��_����gA���?��$���&i��/�B{"xԗ�Tn�}D@�(�&;�� vY����L�m�JD�B�E�J����V�T9�s<؋�К�K�dwv��3K�B/I��>3�����y��ln�$M����g�-[��W���Ȩi:2��<���5�}>|}��i~n1��%=K�b��z��8�v��Eq���{���4�\�陃�`�
�������c�����?w��>���ǸS�O�%y�z�s_��\�� ���@�۱y��v��9�w_����]p΅g�<���*EG���p��v:��j�ڛ��:�Gy�Bތ�޹h�	=���M�Bw{c��7c�����sc\���ͱ�}�V,v�bv�^ ��S?���L��ç�7��n�7z6��;�=�~6�O�������g�����xs>��F{D��9����'X��������� �Wh�֭k��S�Y�|r��=/:��B�W�'��#����Ճ��4#��G���pd������
�����?�k� 8!:�V�)]=r������߻�sO{ʏ�,����I�H��*�ē.א��������g�����? �0h;׾g�ߏ�c˿^���5���'�z���O����m�k�Y8�<-�K6�V�'.~�\��u�}M O�@��x6�<��9�O^�_���+�q�3��-~��Vv�5�#]�w�#OSw�zz�]�s���~��5���G '�@���#��ݕw_��[��\��5k��� p8Ď���7�Ñ���xkX�/�}Z�n��% p�t����;�v���;�;���]t�E�ȥ瑎�
���x�+����3n�ݑ�/ �t�;6�X�aˆ_���}�S.^��P=��G���w��'���!�~��e�Wg+_s�ȵ� ,�t�m�����ߘ\����}������b��.Z�Ý&��P?2ڏyx�G�O�q� �H�3����|��}�_�����ڵ���X���"����������F:ϲ��=�V��Qs�4t�c]=r��������V������c��b�R���G��c����_���١�ͱ(6
�3�3����� $C���k޶iǦ-���-�?��矶f��Ï8:|�0���\���ҵ��G+ H�@������p�;�����Y���~ړ���׻D�m�w�w������� @�:��{�u��;wn��_�˥k~梳/
��M��U�|m�����,y�5C��	 $K�eݺu3qx�Hu�y_��Kv��O<m�Z�����~ja�k�F��& �<��&K�7�a�;޿�=w��|qoo�P�כ����:�w��|�P �et��pݻw�o�Ν_���O�8c��/8��N�ԕkkoY�d�˜��z:�18t���F�Fθ�޿�i���\xޚ�B�����kU>x����%�]y����$�������qx����K��o_��9瞽����E:� ���+�;m�ڷ�6��2 ��:��P�8��qX=49�kw��S}�yO�_!ԁ����d��]k߻�];*�� ���������'._������]�ۿ�_�'̢�w���?���׾5 �V:�<�1z�{��+o���GN���g>�kq�"�̛�0/���.y�뇆� ڎ@�'��x#���^�ƶo�~���7\p��Kz�u�q[�譟Z\�ً�\�Za��:�<;�o������}�=˺�(ԁ��;�[_�ü_�t
�p�\z饳q���;w��ڭ_��╋.��l�<�E�E3k��~�����C�x�Ct����??w�{���]�j��9����>����Ƣ鵅S?�㫞�K��3	t���Щ�oknלּ���z��8�����йB�C�v��Ī��_;�� J�,�k�׼�R���=�o�{�]a���郧�B�:t�B��`c�۫z�su��?�{� �p`�����/L�����%k��9���
� �����X��������}��/ 8�@H@O���ׄ�;g�7���г�7�yڙaq�� ���3��dk�0�s�/n-�� �at���bX=�*�{C���w�����3N	�,_���%˳�tv`����_�i�e�/�t�D-͖��`��<n_�г�7��������t�6z�+��^ճ�׫�~y��M �@H\����W�����/��K�/�������cꐊ�Mߖ��XU�_x�7^z饳 ��@hY���a0�=!ܳ?��z ,�����X=�������O�^u�di���{�� <�u�ך�)aM�)aw�'�U�+|7�/�3��D+���`X~�`����ӵ� ����eKò�C#�aW|�5}w��lW��0_�n���߳�{�sK���Q]_�w��]�<� m�y쪰2��Yf��po�;យ{��=���8>ͻ<��}�W�a��wԮ�}# �	$��P1/�Ӌ��m�랙o������C�:<�,�7XQXq{_X�yǻv�U ��D���E�u^���pn�)�ý3��m��{�N��Nw�H��l�7�������? `t����
gϘ�f��۳�����v������Ŭ�/m�Y�-����� X`�C5�V�̹-��p���s׭��v����n�w__v�(���I_����= "���C�)��ᔞ�!��'�ߙ�N��Ʈ�`�A7��%5O]_�Xr`Y���,�^���zΩ �(��ɲ,,Kò��s�����w�c��]�@�7��'t��7�w-͖޼���7�._��� �����ʻ��2��^9��/<?�����	������y�l�ށ�ү��\35��� Z�@���_��Ϟ;���CaW���+ <7ׯs"u�]ai˲e���&�9����/� �t ����}y_��~f8c.��
4v�E{�Z���s���j��Z�XԌ�0X���aq|rw�T�2 @� ̛fP�a/�`�9s�����} F�����f�e����g��|�@��faE�������� �St N�ft�R<en��|K�\���+^r�1����>��ƃ�=�u�o6���'�K�kYai�aYqiX�X��� �K�p�m���8|���Ν;�o�}��y��]�v��e��f�����VVȲЛ��_�׎��_�����  O���֭[׼�܇m?����{�s�[6�T��f������.ٞ�bV��E�/�x_�/,-���-�Ǐ ��: �z�[��oqxߡ��<�����<8�����=��.L��d3E�~b4C�'���E��Z\XC|`���
]��N�X�c&�h9�����C��~�/����gg^ppf����gN����P_<�8�;�5[��w8]1���ߏ�lQXRX�dK�?/.	]��G�F܊�&�h+�_�=�?=�=���=��C^P�ן9ݘ}R=L�����0�Wo�,���=�a��^�Y^h���5���sa�sī�phk����Sh�zB!/<��q 8�: g�7&�5������nذ8�;?����������3�~�L��j6�/o䍾P�{g�=y1m�1g������Bb���sc�1W�͏�� 4�K��'p=�Y��(��,���y�P���5�f�V�*t�;�U���݅�}py6𪮬;ď��!=~<ŹHL��� �v: <�m�n���mIںu��F�񪹝<����s h)    �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �    h9y�� �f: �r�,�T*}�r��  mB� -�P(\�[ �	� ��F��� �h# hIY��*� �&: Ъ�^�V�_*�� �t �e�y>�@[� @�ʲ���5 @�� ����z^(B���za*���X� �0� -.�LOOO�T1̟_���� ��: ���K�<p�@�dy�oߺu��6n���  -J�@��������Y:T��W����^��s�; �J�@��W�������b��<��eq�# @� ��<�/jG�![c�ճ�hE �@��;�pA�pq��<����۟y�W|' @� ��)n/
4#��z��'ccc/( @�� �b��S��7��;00pC��W7�� �: ����vI��ŵy�;��
: �����ۻ��?�M�j�_�xe ��	t h�7o~�R�ܕeٙ���7c��T*�N ��	t h�=no	��<ϯ��j�2 @�: ��,�>�ÊkSl4T�V{J��G $H�@��)n��?��y��R���� H�@�6Q*��V����<�C���Z-�> @B: �����*�š��?#=�t R"���|,n�<��G�+�J�\.�A �t h#16�)F�Wb�>'�X����~�Z]Y*�� �@�6��������š#}����減 X  �̒%K�h���[cl���h�V;ull�m����  @�@�Y�~��J����3яכ����7 p�	t hC�b��h4~9x&���������HU��= N"� mh�ƍ�W��O���맦��??11�s���� 8I: ������*
�<t#4�C\�/�799y����W � ����譕J��8}Y��8�P(�M�Z��R�tc �L�@˲췃@"��g1�%F�G �@ �X�ʛc\�I��&�x��y���J���r�� N� m�^�_�����8]x\]�?V�V�X� �g �ܦM��aY��+O�[���s�����<���&��dY���\�8�xB��xff�[�l�dӦMw �' :�����J�R��O��Ӻ�������r�� �� "��W����?�ggY�Ÿ��,�J_ �	t �,��<���k�aE\Ͽ�T*����  O�@�R*��V�o��O�E�e�1�?^��.� �q� �ab��Y��?��7�E��b���u=7��  ��@�T,/���}a���O��J�߾}����7 � hÆ߫�j��h4��y�v`����l```���؛b�� #� jxx��J�R��k��c�b��Q�p�: t�r���Z�>;��D���;w�|úu�f <� .���Ȳ�qzQ`��n�޽����^;44t0 ��� ������j��1ԿC}y`�]233��� �x4 h>z훕J�5qzc�z�����7�����5� <� �)�˟����,�~/0�⺾�����1��#� x8 ���#����.����<��8� A� ?d߾}�����'�[k���8n p� ����וJ�Y��w�8��V���J�� �� ����k����y��q�?N��W*�]q�?  t ��xi�X�b�=7p"옜�����ȧ O� �htt���/.
�H?50��,+��c�J�g���� :�@ ���ȿT�՗�y�����mI\�?ݶm�s7l����%���T*��qbb��.�wW�۩�z�/��ꪟؼy���$��c2::z����%�B�Ƹ;�WY�=����O���^244t0 �q: p�FFF�\�V_��	"�Dx����������#���R*�n�����,�>�����k�˕J�o���u��"���622�������"���>11q���� C� �K�\�|��`1қG��&�gw�P�d�Z}V�T�+ �: ��H���/�������&�皸��{����C��'��'���Z��3�F�fT�M\�h^��� @�� �6<<|����='���|zs�R�B�\�� @[� ����1$��eY�9��M\����722�� @�� ��)��w�j��5���ݟ�/��z~lll�ٮGh_ �W��û*��K���q������~�����8}{ �-	t `ޕ�����^�������̗_�V�]*�> h; 8!��ǧc��R����H
̋<ϯ�������ȿ ڊ@ N��8\Q�V��r[�,���%\�?��~��K/� �� �p�Ri�V�=#���0_<qϽ�;��c- �6� 8)�����T*��'�,[x�޿u���lܸ�� @[� �IS.�?]��~&���wW�,�z���;w�|κu�f -O� '����W�n����w�<�ػwo9��9 ��: p�5O˞��x^�XlF���[��W�j�O� hi X�����ر�'8��{I�qi��޼�����s�5�%���~��}7�pë���q���׳���~5� �,� ,�C����j��M�J��m�T*�*��� �$� $�g�7���K���vq�� @K� @2=+��8�/18��כk���q�G ��t  )�r�s[�n}~�����{V��5/��|�Ν;���� �G� �i>��V�=����؜?8�޽��8n �� $ixx�ߦ��^033�ɸ���1+
�ٶmۇ7l�� @�� @��������]��߿#˲u�c��^�o��h �et  i����8�z�R�V���c���fו��; -A� -!��D�{��a���x,������) �: �2b�drr��1��8�U\�7LLLl�5 �<� �������j��y�|����)�ū��� @�: �r���oٶm�O�����,;=�h^R�V�W*�n $M� -iÆ�#���"�I�G��y�� $M� -+F��NNN�d����+���U��g�J� $K� -mdd�ޫ��ꧺ���"��s��Q�� �%����y��&&&^R(���������[�^�q��� I� @[�#��1�?c�y��fgg��7 �$���ь������������?*��/lٲedӦMw �#���244�'F�˺���7���G�*�o����t ��lڴiw�����l�e��ק���?44t0 �� ��C���������s�,[=33Ӽ��G I� @�jFz�V{Y���=�>=p�eA�$G� mmxxx����K�����e����nݺ�?mܸ�� �� @���V�]������)�0;;��8t��t �#�����
�����B�˲�ұ�����ǧ I� @��z�V{M������������i? H�@ :������T*o	߿IZ!t�7��� t�r����Y�]:X��_�e˖eͻ� �@ :R�����yq::עb���8~$ ��: б���;200�8�$t����� t������������q�?��e�O�ر����� J� mttto�Rye��cuU�<=������fq N� �\.�Z��R��E��;��l� N� D�R��J���Y���?� �@ 8d߾}�������/��܉��GGG�g `�t �C�7����z����W��i��dY�<�]�, � p��������[�<�1Fk:D�P��8l ,� p�R�tS�R�.N/"��g �@ x���xQ�^:@�ek�l�rƦM�� ,� �0���������_�S��³� ��@ x###_�V���_�P��I `At �G�e�H��xeW�6�:t��%� ����j���8�`hsY�=# �`: �c8묳���;���������j��� �t �1\z饳�J�q�����<?7`t �cP*�>Y��6���C˲�8�C ��  � �k^�T������A`t �c���s���t����.��@ 8FCCC+��G�ڔ#� G� �,�>�8���7 X �8�V������� X �84oW�V?�o�I�,� p��<���m��s ,��@fgg����j�/�I�P�F��pOh_��,��@6mڴ;���eY�z��zw��ٽnݺ� �I%� �S�T�9���yw��ѿw�������o��@ �\ �E�_�~���y6o� 8�:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $����$%Gy>*    IEND�B`�PK
     `_[	^�G�  �  /   images/9ba3df0f-d630-43f7-8169-617793654d93.png�PNG

   IHDR   d   }   T;�   	pHYs     ��  sIDATx��	��yǿ�sfvv�ОZd����XĎ�;N�g[(���p:�w 
`'X�B�1�������#��:@ ����c��9��|_Ϭ4ZV�EB=5��������]������Z�JU ��
D0U��*�T"��@S�`�LU ��
D0U��*�T"��@S�`�LU ��
D0U��O]�f���� 8��S*V���F���!�=�J��@?��)�������w��ςfܤ��%�c"�4�w�������|~R�o�p9����ƽP	Ȣ'���y�q/����;	+��j�����ܬ	K?��`Bq�� ���}�|a��Ȗ/�p��W��i�>YB���E�h4�nmlj�'��<7���M�ŏSV<��G�Y^�O	
�YNg|.~xE���#�5X����0�~n!�����AD	�o����9t'{@���S�v^��G�1Y���eC���#<����g�����)��>���=n�lX��"!���@=��A����R�󼻗�E,Ə�Xl,�X�� Z��JG�C�����F�o{�#3�e�u �������ֲ݀cG]wh�|],(er�Ӌ��M�}��/�}7ƅ��#�
�Vl?�E���ɍ�:�������lu,�reI�p���,i˵�OK��DKy@ K)�eO^9%[���:_��
#e��>^��?��� B��N>��ke,RW[Wbb�D��=�~D�b"�����;��N��*����Y��
+���a(������ ���j����gƷ�ho��l+�2���%y���l0On�k�7���xRKJgM8���f��n�z3�$�*�riC��u[v`����=ʭ� Y�fq�-����ƹ��2|>�i�>��+��
�j�.����dw��
ZɎ��;��v6LҦ�N�k��(��4�X\�K��|=���ZR�^l_�0�-e�6Ct�Ȳ'�AF͇֡z�El��-(��S[N�u�vQ��Fˀ�s�n{5Gq[O���n�{����g'�U�P�kB����;^�c�� ���|�����;�*�P�W^�9ʶ�$ M��� Ŝ�*lR�$}z��8Y�P�]�5jB�������0@s���D�\ܾ�>o���;���:cg|MVY]�N�V�����h��I�.�-^KE���v��P����r"�*�!ޠ�l��m��S�܏�|�-/��g��������9��Zb�<eh3�t��+��֒[�f	�7�|Ic�@=�z����JZ�|(������=t-�C�~��ֆ=M
ڇsY�E��������`]��LE!�����PNE
���0v���X�!�NI�H06��dmؽѤ����(��a���O���1��~+R ���i쭉��
}Ra��q�:+�G�"3�m��޸�mK��n�cyh��`Z.n�@w�梧��}���m��^�º7v�ɟ�oy��!���S0��܊�������1�A��N �ϣ�z�K�	��s`�O�
=�V�ͩ����RwEV�u`�CA�p	�(t[0Ǖ]H8q(�"��*X��j?�7���q�F��QEր-�`gf�C` :��'%�DƲ�Hd@�?����(�
L�FKJX�����i?BQ>��3����l��,H�5��*L�TIe�����0�9� 3iN��DBwʺ�L��F���>��Y@�J��Ѝ�%��d�NʨȀP@W=� �R͜C���S�"�C�Y˕���R�`���x�$(�0o?l��X��N��;%�u5Vܷ�)4pB8�VwG���B�B�T<��A�kyI�h$
��vʵܸ$K~�9Ս�*��ɶ협1t3c�y��Z��sT��$I�U�	,1�ൌMb�6�V^H�]�c��"��D_q_��Y),���<��u\��<Y����?�ӌR�a'���AH ����%�����D/�$kpL'a����A
�ш``�ɮi���`���/���O��� ���lL��8ʵ]=��7cs�U���>�Xڲ,	�SL�X�V3��TI0H��A�4)�A�ف���P�(�8U:���R����4O�.������@���stS�讜p�R���~N�C a���}� �1TS	�� C
a����s�3˴�X"��Uv=׃���5���^��UV �uϕ8r�-&3�5�|K�1,��C�ـ�M���ޡ���S�zl�Q0�@MM�-�i!'����H��^���2���D���
�V�⺮$�Cs7P$E6A��᬴Q�P�@��_G;�ԁ���x1����ZMm���Y8�8������6&��iy�VY�Pm���]8T?	��2�d	����oC��y3r�JP�@Ё��j���/l��\x�E�۟��)��g����Wbeo��R۲�XL��r<��mnز ���bю����x�TtU�p��Vn�k9����凶�0��M��c�1M:��)�u�m��sgI�e��?�D������d�df_|`.>�:��a�w���8"B�i�f�3�K�\��?���R��Xp.�W�|	a|'�Èn\��C2U�l@PA@�K�(�i�6\���y�I$�Ӱ`����c��ޒ�(h,��M{�vWmd��qa����ވ�K�2Y��,g�i�1�塐��C~G	�RG�pe�Rd@�����EX�/�H�<��b,\������,�rP�`�A�.����0s�#������!*E�ʛ@)�k;���A��n�Ƒ�W]}}�0���.�L�2,�G�����G�i:D�%)���[ x�*��UEWt
��ذ��.Y��O���(�G
d�;A�(ad�5)�.+
�3o�=���[G�#!�����X"B��ѐN�ǰ�X�! �������u`����oow[ Ƣ�y�v.�<�j�^���!(�Ԝ�Q�����!��B
���*�`Bt3ܢ�\t�p���x-t�t2��:��K�E�1���C}�u̇`H��y���&A�Gv\�Q҃�pBm+��<���->�sC�GGa���AD���\O��gR�?�\pUd?�қۂVx����"�\D���R���m_3�Ϟ:���p\o,�;LV���'ue����$��5*�D>�K� �`��
��K�8i�{�b>�3y6�������)�;��l¸	��[2�Z�ף~%Z�/�v.������O�
��y���t�b;{v&<���4f�!�Ӻ� s�	����q�6�0�P֨��ul��Y���7���~���[a执��T�ڤ5՞9��DO��A03���
g(@�s��nA4Pb��Mz������ښl�u�vēj���_o�|���)�n�Ӽ�u<uc��aYx���nߒ��!\��^}/��ϦT�;g�ɭ��ֶu��ͩf8�����]�L�0]��`r�P2v�3<�w|'\���T$�������0�Hh5P�Po`)���*?m�a]�:���{��
(���hgY�$��5�Utk��b�����6�UAׅn)�!O�9�}���Aظ�mxi��ɂ����7��q�qjKc�J�HhQ�a�<�(��h�Sr<i{�Î��|_f_��?Qu������w�݁��&�������}��S�)�ųϹ�˻[Ͻ[���
D� L��4زwd�,�w�oc��'c�6�YBK0]�hŸ����`9&�<62�5�`8F�n#Y���~��TXs�������ƣ7<�Pd@�\~'\�����`#<��0��y��_O%S��;�*��Н���h&U1����r����h��X��s_�-�"@Vd<�O�~�t\+�������l�����Q(�"�߿����۞����Bx��o|�G+?����<���i�6ih���J
��я�acyL��(磓�7��7?�TY��z��Bz` &�8	�r�7}t?���l}����lk�Y������Q��=�vc#�Y���9�o$���� 	������%����*ҷ>����!�u����>��,gH�`�>�y�ǫ�?,��Z�F�� l>�-�	lA�<�^tf����0#��|ӏ@�}��m�����x�� ��a��O��@ ��&�v��0ض��.��	Xݴ�S���Dcz��$l)A��!ɒP˒���d߱�?��ҙ�,x�} u2���Tv #)(�kL�L������̻������0_�D�m�6��L���@���.����1����BK	09����A�T߽�@d		�T�~�9��$O�t0I� LʒMফ�`�|������a����o1�~*A�)Փ7>�����ܨ�)l�UQ@�?�
D0�@ȕ�-7rm˗/�u� �0��)꼺�����/@�X�B�N�
,�a	'x���PW#c�����F؄\�cXh��7����t�RM��n�;�K��a3:χ��a���p�hU��uPG$j7�+��=�����r+��}U<�e˖�[�`�+,��'�`����!��A�x $��(4���x�C����G�z�q�4������y��S�_��L,Y���B���yXh��H3nN�Bͬ;DZ���B�~���X^�2Ҙ�+��B��+W��k��ʭ�i�MX.��+����&�W�<.����P��xn�0(o`�ˏGؔ,�qD��B>Q��͖���J��[z��*|:��
]����@�A��.��1��;p�3�����i��װԖ�_:�}	�����)a%�c�,_.V��hHUT"��@S�`�LU ��
D0U��*�T"��@S�`�LU ��
D0U���W�cfrJ�    IEND�B`�PK
     `_[�e�e�  �  /   images/3d0a314b-f708-4b2c-819f-35c414b123ec.png�PNG

   IHDR  �  �   )��   	pHYs     ��  ��IDATx���	���}����tH��$s�F��`.� �v�aBf'�O��ēd���`q��$��Ɍ3;;�M2�0�F�@�!��!�9BWKBg�������[���V���<�t!d�<���[����l    �8�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   � ��c����Je^�V�ӨՎ�4�����T�ޓN����I�j�S�F����T�֛�Z��ߓK�7��r#�*'�k��p�K!��6����!�5�H5��S�dv�����J��յ��5k� h �Fޙr��|�~b�RY��V��V*s2���T���fh�����K/����sJ�L�X�fG>2��J.����n)�ӯ׳ٗ�s漺�O�� ��	t :ֳ7��[ڿ��B�zN�Z=&W��k~����{饾�oI�ȥ��B�s.�Ri����E?�6m�|��C�|~o9�����R:�������G�ԉ_�B)  G�@�#<�|�	S��s2��ݥ�)�Ri~����
�z&��z=���<zBX�#o�������W*�����\������N?����7� 0a: m��U�Nɕ�Ww����/4?�޼��nE�V3�������3����/�x���7.�x`,��B���t��K���  ��@K[��O��;w~�06vy��؇zFFNȽ�ڔ����V�z�����~e����=wd����������7uw?|��5�  ���ʧ?]|��k�1~y��ة]O>yt�V��]�\�\.�9y��d����fK�]r�c����r_�����`��N��o\{��Ӫ��=�×�=��IS��hq���I��'%�Y!|��c.��������e�k.��W p�: �y��??::�dR���gt���M��j4�OT�tɶ�du=y��S[�;o�p_�����{�;�.���� Da�7����w㤑�kz^y�t���m�@+zk���k���֭���|�������}�-# ��#fݒ%��J�>>ytt��_<��G9������}�$�����f�%�l�2宝���X��b �@`�={㍽�={�?�;v�e�[�i�7����<�d��y��˞�鹧�����֬) �P�qw[���0ix����?�J9?��VS��]�<j�쯿r���4c��E��� ��t ���˗�0�R��i7.ΕJ�&�J��Oݳ�����~w�ԩ_ߗ��ɥk�n �: ����򱱏Oڿ���[����t�w)W,N�],^?+����K/�ށ�So9�C�J��� ڔ@�xbժ{GG�ɴ���J���T��y��?ع�7^���
�岻�� ��t ޗ�+V��>8����^;����*g���iɪ��t��^v�3{�L�O���_3 @�� �k�6�����h����[��M�L�z=��`���ƅn�3u������w Z�@��=��?�wh�fn���p�#�gx���㦭{����.^|gc֬�x�-��W��$����q���*?3mÆ�ɤ� �)��Ξ;:�����7�x�U�N����c{ �"�xG�\��ģ��~{���%ۊD.S.��ܹse}Ϟ��P�oߤI�w�w� �t ~��Wϟ28����L��~V�r��j���Mߵk�����o�N���B��y��=�������}v�o,M'@�K����v-n~]_��UWݿ���sW�y�  � �V��1wt��gnذ�� m&���l}��o�5/\s�ݛ���[v�}C ""�:س7�؛۹���6]+���r�{����O��=�d�-/M����׬� ��@�PO/]��_~���ccSt�\��7g۶_��ۻ��e���u� �� �ѥK�������l�z\��522縑��{�%�|j�QG}���o. �"�:D2 n��=�?}۶�B��
����{��/]qŷ��:���z��  L���W>�����/����w�~�z=3}׮�'>��ŋ������|: I����˗��>�Ŀ�Z,N�!ɖ�}s>5upp��U�~}ѝw> `t�6���ճg����Ӷl��a;;�'�##8f�����+�x�4oޯ�}�-# Ƒ@h3�t�9�7�j2�����^O�صkqyh�ѧ�/���s�W ���&Y�jἽ{��o��3pX�K���m���W.��cCs��+C� ��5n�)���O~f֦M��T�]�q��{�\4���o<�t��s��- �a$�Z�c+W����_��9CC�`Bd���l���.�l����i�wl pt�������͛?�qu�Sj֬L������k�;j�Z5��L޻������^���<wݺ�
 �>	t����fN��S6o>7��0:Z�_tQWH�R�^o4����|���ju`��ؽ����d��c�n��KW\q�L�_,~���x�:@y|ٲ��6l������ �Icd�����LɄt:��>=�m>��'���o(��P��7o�V7n�&�7�C����v]������U���{�x�:@x��?�޷��3�n�.�לq����@;������|�?���8p�Vk���b��zSatt�����s�\s�^xS�曽���"�"���ۺ���>:�8�o�V���?�ߛ�4)�=��QH���w�U7l�T_y�Ҍ����t����}�Ͽ���|k��z�=�� �	t��%���l��+�Z-`�����N��s�f����K�{��*�X���r��gO��z���	�ſ~rŊ����k� p:@���S���d�-�4lig���7FG멞�����$���睗	��U߽�V{��r��;re=W.��e�~�k�r�׾��  ?�@���Wϟ���e���B{�H�;��i���HϜ�i>�s\Еl��|���ꫯVB��9_��zz���׿z�e�=��Y3 �t��<�bŕ�l��Rir�	���/Xp����T*=~��|�?�Fm��J���M���r}۔�{?�56���?��_<��۟ �6:@$�[��Wfo��ϓ!S���֭�����*RٓO�'�ܞ=���ϗ*/�P	�jۗzat��y��~���K?���{� ��xp�={㍽}[����[�p��|�֨T�\nB��g���/��'w�E��K/�+�ח����L��u̶m������Щ]�YW���	t�#���L۸��CC�8����ع���?BoH��ܙgrg��OΪ��}�\{�J�no4R�v��Ć�:iݒ%?���� �p�<�r���7m��\�8=@$�C��@���Ϊw5�]�j���;8T�MC}���g�V����+n�t�����'���Ǘ-[~�֭�W�\���{��0KϚ�),[֛�S�|�;����_NV��M�����V���+~��k�
 t4�0��]����l��k���d�P�7B:=!����z��{�\PHΨW_x�ܨ�B;ɗJSl��W�W��7�֮�3 б�8�@�]s���ٺ����(�~B�ܨ��]KϞ�k�ԤI��G?ړ[��P~��R�����=w��-��;�����O���_�v�B>�{��O۾�� ��m�]��@�W��=�P~≱��/WB�H�뙣�o��/^u��S���_ t�(������Sz�o�J���	Z@2I=�uV!D,5}z��tio�3*�G�������Fj�Ν+_��)']z���6��"���߬\9u����CC��Z�-����O~2[}�����ط�-�v��]�ox��5/���p��5� @G� ���իg�߱���������H�18XKM��	� �Je.�g�;.Wy��R����a�ܔ�{�
a�+����'~�� @�� ���eˎ=f`����QZP2�=�*���L*w�]�Nȕ~�X}����	�N&��{ցg���go��cg�r�H ��	t���[˗/8n��/7�|V�u��)��CJM��)\w]_�7*�*6��Zz������ү�~��V}��;�� h[�0z���N�?0���^� -�>0���ɖ����|���c��|�����{8�F�GW����w��f �-	t����+>|��m�+�����޽���h=�ӓ-,�˥�_ܝ=��|�k_���ٲ��3<|�����z����Y�- �v:�a���U��ݶ�ϲ�6�܇�]�����3fd�����Շ�u���=z��>�߿��5kv ڊ@x��X���9[�~)[*M�F�۷W���.�"�9������7�l�JO�O6��|����.Z�fo �mt���[+V3o`��\�4%t�Tww�Q,6m��B����33]��d_r6���S�Po�r���s�<{�י��>:�{��s~������d����rg�](�}�H��7�2��;�y�F��H�q�v���_xaw��>v｣�Z��{���7޸����^���D:@� ���n�9k��;�FF����s��.�NM�t�<ra�Ҟ���<���z=4v��o�m�?&=o^���þ���X{�Jh1���'|0�/������׬) Z�@x����O��i���##�B�K�<������@+�]+V�6#=�J������@-�Ɓ~Pww���Sy��r��(�� �I���׳��y[�?�~͚�����]���{g|����cC�˞tR�Ќ�$���罹O�t7��x�#�x��CS߼�-j�t�����}�T*w晅��ٙ�u�FCC-�E=eϞ��J�Y��? �,�p�7ݔ����y��gK����W^ٓ]��g����>:��䒮�7�9hK��[���r���K�OM��	m,=gN���~�o���Zj���ݻ/�k����}���$��K�>�'3��]�X�Sr��/�I
��Z��Ї��{�ԫ����m*�V~�R��̛�͞yf>{�	�d�ZhG����{���O��F��8jǎ��.]��{�����#��w/�쌁�e�]5���teO;����W\���'����V�&��7��ʝqF>{��l+�T*�]�Y�ҥ��/�r�%*��h����'W�x���k� ���3<�t�����Ц2��e
K���&O~�[�3�Taٲ�◾4�jgwyo����+��ח2'��ϟ{n!�K�Lv��|���̌�u�H�|m�����۶}����.�瞧 -C����Xq�1۶���|��M*r�ߕ?��� ���Iw]{mo1��^���j#�_2�<9�P}��r��=�hQ!={v[��HϘ��ᆾ�=����.�L��ưo�ك˖��rݺM���V?@�GV�Z�`۶���V�Ӷ��S�%Kz��{X��JϚ�I�H/�];�J�v9������R���j%���r���f؆6�J�b[�����C�V�����p߾�z����}�-#��	t����u>k˖�j����LfΜLa��ԤI�Oمs�f�U��m��;Q��H�n�PɞrJ>ᅅ��Z�p�Q����N��W�%��{����n�t�m���ݑ?��c���^����=22/���9�
�\�5�ӷ�m�={jɊj�3%������/��g�]H�S���֟����Ԕ)����z���'����]]����3��	t���#������CIe2!�U��SN����͈)\sMOchh��c�U���Q�<�t���˕��w�N>9�|}��;�|�Cyݺ���1v3w�X��O��v�_ �%����˖]?g��O�6���I�/��|��=?�=��������;��p�|����^�毸��Χ'�9���}'������ڶ�X������� @�:�[�^��y[����_������W��M���{����]�?�+_n�UF�_m۶���x {�y]�E�
�}�b�����v}�}c_��p�oDe��¼;�t}�Ջ֬ DG�4={㍽�6l��L���Dr�Ua��d%�H~�s�����)�w�h��ֶ�o{,&׽xqwj֬�~=r��f���~�H�S D�0::{ڮ]�|�� @tZ�"��ҷm۟��P�ܹ����~��!{�����ݵ���� oi4�&Fo�u8��r���ʫ�i�2=�_�W������`ԑ>iϞ=w�5�s�׾�� @T:��x�oM� ��t:�/��;w���ݞ�aP߷�^{�5���;�z(?�D��ys��dIOjʔ�=���<9���O�׬iE�sv����W�xn�ڵw �!Ё��|�z͜-[~!����ڗ-��.\�1J&�/^�ӌ��Ʈ]��#j۷�F����WvgO<1ί�C�������WLΤ��o����۷�ރ˖=s�u� Q�@����+�6_��A�^o����S]�^ۓ>��\�Xr-U�u���!�S��h�R��n�h}`������V��G�������pĈ�����㇆���M7-N�|s��'@'�@��������C�Kuw�����7�Z@��ص|yO�_I�7Ï�<�l�鵃7L�|Dn x�F�'>�;��/G=8�op������j>u -�b�p{f��_��u������%+u����[j@z��\rV���C� o��曵⭷(,_ޛ�?�%_���z��^3񎑣v��_֯Z�Т;�|$ pD��<���K��8gǎ_-�+t�:T+d�ػ����xIԖ�c8����N�n��H�`�Z������r9�HO���}�x��/?��[F G�@:�m�����K�Z�
-�Ӣ�[2� 9g|p���M� o#�3�����޽��%�t%�C�Iϙ�M��$o6$�>1*���*l���ͧ� 8b:�QNٿ��{���v0���{���e2��%KzFo�-��q���.���z���zZqx\�M?�|yoi��hg/�x�ͫ�����Ϲ��� G�@:ƣK�^q��@hao���%��C���Nw�X�[lFz2�;�;�|������Hr.=� �����G?�]~��Xg/���#���G/Z�f[ `�	t�#��ս�������W��zzRݫV��T�&9�[X���t�]#&���$�!J_��pr�;ys'���g���*�חB���r߬;����k N�a~����bqFhQ�R����ZmZ���=��\㢋�ʏ<2২��Q����dBz����"=��]I�W_}�"4e��3��.ι��� �Ph{�W��d�ƍKC�Juu��>���d�9��ܹ�{�Ԓ��~���ݵ�d%�������T*��暞���pm��(���y���<����k�� L���dj���[��U���2�еbEOz֬���ߵ$\����>88\�2\�G}Ϟ��HOv����T��r�T��z�_��p3ԣ;ב)�{�����O. 0a:��N޿�s����C+J�B~ٲ������I2�T!w�Í��Dz�;Fz>���;����'ׯ������h������gM `Bt�m=~�u��޼��Т�_ޝ]�0:P�����b�V���ص�6v�]#�d�{�MwOϜ�)\uUwiݺ��F����k�o<{��ξ喑 ���@�:j������Zr�9����YgBK������t｣�R��$��J��3����j��gO<1_߾�Vy��&����;����_ Ɲ@�ҳK��Z�m'��|���]pAW�`�$C��O<]���W�=��ha��d�Ah!�K.���U�m�Z���k��G�.���{�}( 0�:�v_�z�Qo��OB�uT&��-�)y�������&��3U_z���4i,��ݡ�$��,�)�z���H\[F����}�~���K�_���F�q$Ё�3m��?�T����ח.\{mo2�9�wޚ�^ۻw89k�g�<�T)=uj:{�i-uL$�|X��w��ۇ�Qb�=22嵐�_i>�| `�t��<�bŅӶl�(��l6սreo�=��7-�������/h��Ƶ�H��=TLO��Iϛ�2�u����R#3kV&���g�����^���qǛ�q�2?� ż}�~7َZL��+�;���(5yr���c_��p�]���kd��G�o�aR�bR�7�����wגG�3$	�F���O�r�g����6��� ���@���ҥ��o����;�B�S:�:�w+=wn6w�U=����J*�oi�ڑ���Kv��O�Vk4�7߬%C��;v��V�>pƞ=W=�bŇ.Z��;��N�m����6mj�k�2��e��́C����h�N�WR�$�ˏ<R�_~y�x�Y����޽�Z�Ɋ��=���v|��9CC�k>[ 8�:�&�����i���z{S���{Z����/������qctWR�ʳϖ�s�d�'�|�v�$��k?�E��k����w�S˖���u�n Vhy.[v����W�V�J��%Kz�����V�N�����/����(��)=�P13wn&5eʻ��P�7##�ڞ=�z�M=yT;}X�={~�����O_�� 8l:����t��R�)��?�+}�ѹ�{W(�˗�o��@htt+q(��F��{G�����q�J��O��љ����6��^ ��@K{|��s�n�z~h!������k�7b��1#�=���Z3��O=U�_pAWG�g�w�a}��Y3 8,:��f�N+]����>�5;٢x_���ʓO�U7m���_3/�X����)S.������� 8,:в�\��ɯ�~fh!�+��N����
Q�V��~�T~��R(�l=�ݩ׃8?|f�޽�U�>��w�	 �ohY3�����-��=��|���w�^5���/WJ�<2��D S�v�IV�- �	t�%=�bŕ�6o>�U�OS�&��]�����uk��������Cdf��}�W���w��f �}�@K����7��X=O�T[��;�:xwJ�z��G�*/�P6��ܢ1����l>�� ��"Ё��~Ŋk&m�|B��Z����]��.U�x�R~��b����!r���Y�~�깋�c{ �=�@˙�o_묞���s^�8d���z��(V_y�������8��ͧ�< �	t��<�|�u��7/-��Lm/Z�̈́T_z�\���)���g���W?�z���ck �=�@K�58�2�3ٓO�e,���PT���=Vy��R ZR�V�MN��& �t�e<�bŇ{7m:)��TWW*�����~�w�J��;R߳�Yshq���fݒ%���w�P �]�@˘=:��C��{��袮TO���?��-�_�z1YA@��T*=h4�e�� �kh	.[v�m��- 3{v&w����;jT*����g�}������_�� xW:��˿�������J��e�u�t�%V���dJ{��Gj;vx�m(W,N_02��ͧ�= ���b�x�y�i�v]Z@��S�|���w�ص�:z�]�ax�yshc3����A��k^Dћ�h�r�\��Z6��_pAW�mU_{�R���Q�͡��8p�˖-9ݺ� �L�Qk�tSz۽��
- w�y�ԤIý��sϕ����m�b���?k~� �@���SO��c��!v}}��9�?��h����b�g��(���?��+N�x�ڗ �D�Q�64�B�_|qW*�3�����*V_xA�C'����J�_j>�L ��t Z��Z�p�ƍ'�ȥf���N:)�;I�?�`����s�`S��r��>�[���JE�C ЁhM���
L����p�U�;�Z�t���8B�\��ٶ����� ��:����3��x��̜9�����@���7Z}�Uq4���䨒@8^TQZ0<����ؔ��v�T��y�^o��[7Z{�5q�P���iɑ�K�� �O%Ё(M�!D.3o^6{�Ξ'��g��9�������O5��z ��@t�q���m�|Z�\���]����㏏�����/n�t�o�n�� xG�Όb�b��=;�=��C�*�?_*?�D) ��|�4��'�\�|z{ �yq	Dg����!r�.(8{B��W��*��a���?��@T�X���ܦM�C��3f�����g�k۶U���7� �L<sݒ%���w�P �m	t *�GG���.Z�������=��4j� p(ҵZnn*����� x[�ʤ���C�R==�܉'v��yr�����6FG-��ʤ��A��#�D�U��ɿ������gB&�ѫ��o~��lo �R߁���ʕS?z�]� ?A���9p�?D,�Ʉ���C���R����NxOҵZv����5��� �O�@7ݔ�瞨��gN>9�������T߽�V���Mlޗ��� �ޖ@���SO-]P*M˝uVǮ�7�����w��jչs�}�<u�7�\t뭻 ?B�Q�:6�����ٙ����=��o��� �>���L~p0��? ~DǾ��qp{�ڵ煈e�<�cW��[�T*/���9p��8�ls� ?F�GܓO?������|>�9�Ď�F����׊�ag;p��8p�7��{�-�� ~H�G\_��4D,w�)�T3�C�<��h��[ہ�*��^ٻ����[ ?$Ё#�wx8���'�ܑ����^�T���J ��Ʈ
�Gt��zt���=��>?D*5mZ:=gN&t�dk{��G�8�>; �#:pD����z�w�gO9%R����^y���訃���)�3[����� �A8�zFF.˝tR.t��޽��sϕ�8�[�� ��"Ё#���N��̛�MM��q��K��F�Q���6it�� �	t��y���?rR�׫e:p����k�ڦM� 0��������<�5� Ё#hZ��,�*�
�:+Ы�F�� $]�����U�_	 t���97D*3wn&5iR����C��gJ��!w���T�"t��:pD��ߟ�~��cB��'��Qw�'תU����	�S,F;�`�	t��)/�]�E��<��v����sϕŢkՀ	�5<<�9t���Q/@�x��˗�H�f�J��w���F�l�8bR�zfZ����{@����],�"�=�����X��w��GTo�|i� 82�GG�He�=6ڭ����s �ccg :0���Ss7Fy�y��+��3�c��W�="�}����M7�S7��&	��	t`��T�W�He�9&2�T��Z���3Vρ#.S�v���n>�N �`�p�b��!R�CT_{���zD��ZM�C�@G��@<���B�2G�1���=W ��;7 t��y!
�!����7g����SS�t����޽�ڶm� ��bqA �p�P}����^O�e�=�c�'V��v��ȏ��|�ӟ.���/��t��y1
ġ���P�Tz������\�Vy��J �H�^ϼ�qc�3���CuċQ ݕ�I!R�y�:b{{�WʡT�|D��VKΡt�c	t`B��ƎJuw�R�'G���p�����s J]�ʩ��	t`Bu���Jϛ��T���������aP��:0a��b�1�M�zB�2s�v�����P���#}`�t`���R�He���@�����@����GW��}�w� :�@&L�T:+�(�
�Y��>�mob�h4R�r9y3��@����*�?"��4)
��g{;�
�����\�t$�L�\�2'D(={vۯ�'j��f{;�|�r\ �P�0ٱ�!B��j��u���@����Q�C	t`B<��ߝ{����m���۫�Z- �.[.� J�"S.����=㙙3���y��9�"�Ҵ С:0!ҕ�)!B�L�o�ĵ�ږ-h	�j��5�S	t`B�k��C��M˄t:ʕ�åQ.7�;w����t�|j�@:�@&D3��e�Mk����ρ��U�����p �0��ryn�P���m���@K�T���$Ё	��Tf��;!�w�|��|��� Ё:0!��r�Sy�0 ��{�@ZJ�\� :�@��m�����/�����Ɓ�F�� -$[�N H��nA�:;4�MJO�B������g��s���j�(��ow�J%�q==�������a԰�hA�j�; t ���t�e�;�f����h͚b � w�o4QNp}}��v	t�%�FG�7w_ D��.[��Juu����P�7���@*d��$w�t���\�>=D(���ց�m4jЁU��j�8w�z}j�Qww[oqo��s�e����t`�e��(=����+�����t����q$Ёq���'�����Ȉt�ee#=0�:0�R�zW�P:�o�@�@�J7�B:�@�_��1���=�mqZW�� F��.�hdB�R�Bhg���,뛻 �H���q~��f�z=�JVЁ����!Ё��f���#�T�oq��ha�:�q�|���t�[�C&�O�)���-+�u*Ё|��]�g�S����+�Z�@�r�D�zt��J�C۳�ha�Dw�����J�
:в��/O���.�@o����z�ahai�t �����~���^w:���6'�'	t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@ xc�z��h����N��t� h{ ���̮ry֑��q>6�P� h{ ��f2��lv�`�:5 �8�  ?Ŵ\n�Z�gF��I Ƒ@ �f
���R�T�w ' �gH��8�P�5P,U! `t �C��>��k���؜z�  ��@ 8D�T�zT����RiN8�� ��@hc�f@��j��\W:]ʤR�����;�g����k ��ЦJ�z~W�4�B.@�I�Gz�щ�3]��x� m�X.wm/��[pis]�tqv���H�ٮ_�p� m�V��GJ��Z�b�m��N�%�Տ����5 '��&��jn��:@>�.%q�:8j��q� ��@hq�F#526�]�ם5�#4_�T���w%מ��~��E���J����Usg�����)vN���C��5 �ТFK��r�jK-�q�M����HVғ�Ut �+��b��Z&Y5o4� "��d�:�NWB��Q��Y*�� �����˅�JŴh:M2���B:]J���!q�@ �t�P����cc=�F����1;��ՕN�B�!�v�J�Mp�p� �s}�lf.��'�)�%q��T�U�� �)ק���r{�����7K��c�zw ��D�D��it�������p�ԮRiF�^����J�D��it�f�N��B��T*�F���  ��@���� ��t���\n���Je�jur �q �"��4�;��U(���T&U�S ��p�>�V!�����w'Pr�����޺u���־"6!�@�ق��8�$�U,���L��=g�9�%3��ɛ����x&�M���l��xc1#��lf�@hi��[�w���/T�,KH���ߪ��{�$Cw�������C�ðk$ �"��Ev��w�f#8t��mW�zސU;��<�0��Vg
  F�@�q|�;�eUM��Rf�� �&!���8>���&��qn�Db�ry۪����+ �It h�O~'��pn&3�XV(�DQz[�B� ��@���4�������m)�
�@~�t����  4� ��i���yڶ}1PE��JeN$��
 ��#��A�R����ߣf���=ۮ���(�u��� Z�@ � Sځ=��<�8e1���-��@�7�  -C� ��tݝ9�)������R��+�&� ��"� @C��R#��T^T��J�W ��t  �0}��h�뎋��*���(�
   � @Ct��Ā뎉�vT�3JQ�  A� �i�y~���C��@>�  ��  `Zem����j���&��W  0�  ��g��ٞ�C5��=cA�/  �@  �"mە��7d�6G7O>�F�`P  0�  �,���M��bfwT�3  ��  `J�`^&����@�0�U��  ��  ���Q���m�e�b�ry���  G� �Co4��\��@�(r�U*�U�}  �G� �C�t�{�]�Q��Z��!� IB� ��R����ۮ��B��Qmy<  �A� �I��N��9NIG���\�r� H ~x ��6��]�S�8�\*�	D\  �t  pP�S���T*/R"ֶJeV�i  �t  p@q�������(�  	F� �wԝJM��j{�2�EY  �t  �_9�.�tݝb�8��Q�%  �  �SƶK�<oX����Q�#  �	  ���mW�x�v����<#��7} @!� ��o�s=o��8���� �  ��  v�o�y�̐];V�<A�5� @"� @M���r,+�0;��3 �6E�  �D����͵�@T
��P�:Kj_*  �@ ����<m۾�Ei� �	t  :����=ۮ���(Jm�Tf��|  �� @�R����ۮ���(r�T*s#G  � :  j����$
�r�V*s�s @'!� �@��ΞT� ��܎�|v �
  �@ ����R�}�;!R"��s_��  �at  :HO*5>�cb ��*�Y�(� �D� �!�l;?�uG�PC���re �E� ���]��y�b��ʌR� �F� ��<�.���b�a�(DQ�  ��t  �Xڶ+s=oȪ-�6�N���^  :  �*�!_59��|�g<�  ��  �!G$���ٵc��3]#A0(  `7 �6Gy8��9���
a����  ~� @�D"�mb�Rf�W��9  �@� �>T�mA�"�rl˒�R��W�y+��ry۪��R{  �@ �=�l��q���ݶm�+�ű�(��S�]�[#��J��U*�9  �@ �d�h,�T�@�\EV�+���r�ߧG�u�����r��Q��q����  ���  $���q�W��c)�� ��)ǩE�mw��!�o/T��Z�̉j� �wB� �`^M��*5����n�W�������1��1�r{K�<'�~ ���L  *E��*���^���G�-�*��@hY�  ��B� �@n�^�@*��e�G�9  �B� �0)�ʙ(�C�l�/��  �I!� H'�*z�v1T�q�B��  L� @B�QT�EѨ�d۽�ee   �p���yٶ{��
  8d:  ���
rQ4"����S��.߶s  ��@ �`�Ra-Ε22Ϋ����v�  �)#� 0�R���8�#1�oۙ�m�
  �:  R��8�m�B1P`�^ɲ�,  Ӆ@ �0:��ȹ�T 
,+]�qn��  L'  ��8M)勁�8w���oQ�  L;  �d�h<��(��T�8 �at  �ḫTYY�S���,[  @C�  �����R%1����8 ��t  Z̍�B:��b�H�.�qG�#  ��t  Z(E�L��@J�*;NdY�/  ��� �ERJ��Q4.�һ��q�
  h
 ��������綝  �4:  Mǹ��:C��/�,O  @S�  4��T���U[�m������  �t:  Mb)���[VV  @K�  4�RQW�#=Ul�ˏ/  -C� �h��yղ�U��  �R:  �bq���J�b ߶3��  �r:  ��\���(����J��g	  0� @��K)U��.�6q �At   Ec�(����8w����9} �At  �Y:'\��b�вR%�1  F!� �F�(�{J�@�e9E�˲  �@ `��QT��� Rq��  ��@ `�J�2Q4!R"���8�  �"� �"'�*q����t��g �,~� `8~X@�ahEJ�	W�����:C����8w�������D hk: L#��AP���=G)?kz��vZ�h�ue�XLg���� �- ��5��8W��w��:Ȇ�U�En�����	�F�ZM�a�t{��h: �' ������wK�0E��y�qz��ڎ~#P��g=/ȥӌ�@�!�`
��Ӫ�;Q1j�)��jq?��ʶ��[VV��J�JJ�)؝���e�F `�t 8DLi�<���<�C�@e���m�K���M�S��T��7�  �C��!`J{��q�G����V\����8݂��gJLy�6A��$0��c�8M)勁|��Tl�Wб��w=�ޓ�2� �@��Ĕ�Ε���8Ϋb�����m�	:��գ���d2�� 	E��A�@ǹ#�8^��q^��-��w�P�g��H�#=�F�  �? ���+�i�Jb�вRE��b�P.�a�]�Ǻt H ����-EyO��(�,�8ǁ����Ql�K�� �`Xo���q�{QT)˲u�K�(��ץ�f�UǶ�t 0� {�q�G�)�T��	1���mƏ���A��Kכ�q^: ��@�=�͉��ޱ]�D��m��8z6�>/=I��ccG�s���;��� @� �`6��lvU�Y�b ��8�#�r��y\�z.�6�(r<��������o��� � : H{ĹU���퍠�e���߀"�o��(2rZ��[Vƶ��V�,0J��H*���3	;�{A`-ܰ���>��n�� m�@���i���mWu���ʶU6����W;�-�<��M�R�tM�𮧽wg2���T�z�'߸��%_��w�
 �1@�R���U��_�z�w1܌��t��G_���+g�������CE��H���8���q�z���\��H��ysߋ?����e m�@�qt��K%��8��g�'!����ү�}����B �� :���8��t:���tJJ��wU?������.�����
 �@Ǩǹ�e� ~_=���t�2�U2֜���?�ɇ�r�M�	 �@G�q>^*��04�� ZLG�~�4}$��Xt�O?��{��r��h':���wk�Mk'����n���s�l�y��{���$ �&t mo�\N�N ��{�\vM?'}�sϝx�y������� � ����L}�) �I��[���<��)�Nɜ����q�����A  �t mKǹ�� �!)W�)�a\.�66һK%g���7�O� �@Ж��M%q SW�TR�e���b�y�7�\���{�y� @�� �N9s}C) �iQ(�]'�t7���P�=��}���W����� H(n`����� ����_[��k�m+1P*������{���&�^�T:����:� ��!�ۯ��l��ץ�h������>?=Y  �t mC�uE��w� ��0�E��g�/|�ٕ�|��]q�-� H@[�;�s�9 4�>�Ro�i���nI�#�|㟯���/]sME  At �ǎ� �\���>ct4=����OW	 $� ��H;�@��9]ǉL�4n�sϭ��������w
 $7� Ko
��T� Z$�kgw1��V�s��#� �@�X�ƐM� �u�����;���@�6o����>t�_�uק �@�H�j���� �Rz�t*ŗ����>��Ǯ�����k��, `8@���"S���J%�r�Ho'��.���/�p_�t� ��t �����r�8 ���F��������Q�x���ꭷ�% `0@�*֝��j��=�C�{����3 F�H}��y� `.}쥗J�&�6��7����/�{�M �P:��`j; ��ԣ�����O?}U�@�0� ��I�����l���;�5nW������?��5}�]	 �@`<}���M
  ��k�>z��]�g<��'���K��Uƭ� nx�@�@�(�,=ս7�5n�����������~Z �0��0��&�G� �(~��rS�H3���?v�W^�(: �� �)e��U^�  ��;�JU�0���_?����' / c�q�1 $�~7vø��� �at F
�M�� �x�n�Gѯ��?��w��9 Cp��H�J�3�����+9]�g�z��������: ��7 @[�3��4wǶ�E��}{���;����m��� �t �)2� ڎ��ޓ��b���^�j�@�07� ��G�9V �O5���a�q�:vmΦM�x���ꭷ�% �b: �0z �K���mX�;Q$=o����� -ƍ0 c0z �z6��[��������]_]��  �B: c0z ���wg2F�E�V*vjh����O	 �7� ���9 t=�����s��6n�3�#�����@��;��6�>{h���.8�+���) �"�h�0�,�=��a�(���x�6���)��et -�w� @G���q�P2c�Fvr�R:���g�
 �����L��b���y�}�on��j� ���=��� @G�v-orS)��E�n�����@�:���0� :V%�}��7	 ���e��j� �����K%�k�����g�&#���� �H���Qk�3[�|.~ �4��e|F����BM���[�	 � ��%��@l �K����c��LsH}������  �D:���p� `�3!�Nb��qj���?� ��@�Lo ��YU�N�I��m;^ ��t M��v ���4�H)ˤ��������/�����# MB�h�*�� �������V��7���~Y �It MWe�9 `/&���� @� �J����v ���4w��X�9?"r۷/ h"@S�9 `t���T$��߹3��W\�}�k* M@�h��N�  �E�+bL����Ro����� h@S�͗  �&����� ��@�4�ctX ��[ˌ�! �$:��	�s ��ah٩�9�>:�# �$:��a�9 �@L[�ޛϻ��zu�W׮- 4��iX 8����>RQ$n�pq��� F�h
}�-�� ����s!�4��)BF� A���7���cc�
 4��)�  p��Fqb�t�0  �:��	t �A���k��c���3 M@�h
�6� ���,�q�]��� �� Ma�zB ����+ˠ@�|����|�]_Z��y�"�4;� �~Sל<�*΍t E�h8F� ����5-�S��) F�h8F� �e�ώRi� @�� �t �d����*� �@�p� �$���$��� F�h�0	t �����S.g �@�p�b 09ƍ�W�i�#�  `�ݭV]�#�4\|��: `RL���\@� δQ  &ˊ82@��   0�io�::�& �4\��pW H2F�4�   �E �F�@�8�DJ���|VmO% ͔��R�?��T HČ�h@��x;�&e۾ hk�(4D��M{��`t��1 �G�h8}�e�] �x�&Ёt ��M `Rt ��@�p��a��� `��g�Q�nY�_ ��t �( `����� ��, �!�g��C�h8�v� �Oq�8�D�h�0�t ���o�_b֠h@��7Y�pc ���7wt @�: `��04*�A�:�����tZ  8Xq�S� :���|�FA  ��Ȩ@g@3� �M�  �p�
�C���ᘦ ��H��0��t Mዸn� �wV	CWC�h@S�J�]�"� �!�� :/~ ����k܀ �@��g���s �bԋ��U��"� ����@�,:���;� (qL<bM	 4��)�Nm�6� `ߪQ��� ��@�4z�8ϲ� �~�?+�[�w �B�h�J�=�!� �U�V�?бx�4�M�ۛ�
  �cZ�3z���z���.Ge��V��| �?P�2�G���t M�o�|�tZ�"  ����ƶ9�@�� ���^�qt �(��h:��*V�i֡ �E/��� ��@�T�j�f: `o��?7�kОt M�op*Je2�U  v)�~F���sF�4�����j&�y: `�|���� ��@�t�rٝ�yLs ��>� 0���s �@�h:�� �T�}�v%����%�� �3qz;�h@K�i�3=O  ����q��5F����%�4��RY��@g+A"��s��f ���D��e�; t��r9��Q�:��ɗJ���c+
 �㔢(��q���s �B�h�|t�:θ  :�x���0R��t -5V,z�== �,A|Z�T1�� Z�@�Rzj#��@���~��@�J:���S3�� d�T2ns8��h5@��e'�fݔR�  �^!���(2��g�3�9f@3� �0Z.w��� ���Rɸ��5F��������y�Tm�  @�*FQ����-�>��s�f@�� �1����;* ��5Z*w���N��5��q ��@`��b1�����J� h;�(ʚ8z~0S�#��h�1�<��jw��	 �팖�F�v�����h�QF�E���߶�� �6*Je�ժq���������% G�0�E�V{Y� �eg��-�rmy�N� �@`��B!�30��� �&��禎����X�J�?
��#�ig��3;��) �DS"��B�ȝ����̞N�1��#��P.�*���,�, ����� ���`Gϵ�u+ F�0�p��=���@��
�)3b {��G�̸ @�� �������l�  ���Tz��&���zˮ 4��h��|.��W��5 H���7Q*�b�Ɏ�ka&�U ��t F��.��fzވ  cG��#�:�@�L�e�#�O�����l 	1���z��HǹeM~�:;��_ ��t ���P�Y��SS3 j|�ԍ�ɮ=ע8�+��� �@�~X#�j߀�
 �X;��>S�K=���J.~�[�*
 4� 1F�t����*�Y� `��0�)W�FNm�e�\+wuU ��@�(C�|��������3 С�����|Vu�q�����)t �R�}k���� �1yj���P��k~O�F�& �$������e-��� `���oǩ�uaOϣ M@�H�����E}}[�P  -S���~�T�G��X�=E��- M@�H�(�d[�00/��! ��E���|�l����l6���� h@b��c�t__*5& ���Q*��Q4����q>�����`^�xC �t ��3��f~������%d�; 4�X�+��O7�T7���Θ� @�� -�h�Ȋ]9����[ @Õ���7H�`S��^����A��!�$Z�)��>�'8�؞��hX~�ɪ  F�w�m|��u�z�|�S�5�7��Z �It ��J��GמGQd٧������x��� � Qܾ���~S�;�t�O��y���z�w�� @�� �������!� ����g���׏D##�  ��P�4�����i��ZqΜ-��K �B�H$'������߯�v*w�y����Ǣ|��! H���j�R���k4]S��*3f�' �D:�D�]�R�tz�wae���;�{�[�R�� 0E�a�3V,��`�9�]�������* �D:�ı����Nz���ݝ���GT�{��+� ��)DQ���DV7�q�+�^w�� MD�H��w�KR==��X���>[ K�`�*Je��ǻ�p:Χsj�V�;w���� @3� �ժ���R��hQW�>���  ZU��2>�+�����5ݪ3f�- �d:�D�-Y"ޜ9=L��_�.]���z��+ 8 }��汱>��SӦ{�y]�J���� 4� Q�O9e�������c{��ձ�/Y �~E��l�7=εFĹ6�`�ȧ��z� @�� #=c��8��� l���ra8V�կ�t ؇ �7�:11���g�k�Xw^W^��'��c �F�H=znM�n��};u�I}�(+=�4[��j#�q��A`|�7jݹ����{{�V �t ���r�s�qS�8z$=�jU_�q� P�Gη��'b�Q����,�5o	 � � �N:Ilם�G�re_��$ ��j����DĹ�J5����p�ϙ��Ut Ƴ⛱��+��c�H/s��\Q �C��ڷNL��oGE��_ h��z�/�TW״�<������l�dY����4
,�ջ�')��)\�؂c�^wݛ -B�0[|3ֿjU�>��H���re۲"�PQ*�el�7	G�i�ܱ}O�E�n�� h����^q�9�9��B&��cۡ @+)��6>ޝ�8o��{*�r��+V���v� @�� �揍ɖ�fi�y�)�q6|ߨ��]]��m mh<{�'&���ޱ}O#G�_uUY ��t W��}�x��e���\���9���ם�Y��pN:���yo�I���.�?Wy��/ ����j�a(S�N��%�����s�mx���t.��<׭
 $\��kW*���+	��8�F.�˛n�G ��t M�o�� �Z����l�?Μ��^,�� �L�� +�,g[�0P�V��{53ε�ᇯ�'� h5@�LG�O<��D������Pv*��H���G�>+�c� $�oY����ޤ�V��8/wwK�/���V�V#�4���#}*jkҿ��ښt�uz�wx+��� I
QԵ}b�+);��5��uԯ������t MU_W8�H�Uټ~����ǔ�N7�n���{.��Y��tcAз3��$aZ���ܹ� A�h����o��[n�yq�;�L������0���.�q"{�T,U*�Zo��"ε�c�y���A �:����HߴI6�]+�?�q���6��R��֥wg�e۲��8 �F�2C�|O�֛k���(�R�/ 0��e�+ҫ;vȦ5kd�(oΜ�����X>���媜��Ւv���Z�ڎ��~���L � :����H�yy��k�ݳ6�nO����S���>Bm�XH�v��q9�-�L �0:���7h��N���\��n�If�}��]��)w}zʻz�;��h��R٭cc=Iۥ���q�y��׭�O �0: cL�9�*����y����f������w��(6vy��5��}��BZ��q�l[£���<�� �it F��H��eٰA��Q�s�9?+�N����y���3��Z �U���^?��V_��jÇ����~�N ��U �2-�˿��2�#Q�������o��~��t �E����~�H������L��0�RGu�l�  `�ֿR�>��0���)}��[oɛ�]'s�H�.XдQ'=�^�+��p�C�[��mb"���)q��8�g�r��{ eƫ% ��8�ǩFzm��u�d�=�Q���ִ�� l}�� &�F�5۶w���Z%��Gq� ��t F�7vz�E��O��#���j�����?�f�K�M0U���B�����5���tS�Xq����� �� ��o�t�O��tm��g��}��=�<�h�hz���l:͹� �@7�H��;Q*��p�����`e�I'}T~�C �� ���Q��Ou�ʶm�u�����c�m�U�Rq*�j�+��]�� bQ�3<1�M��{j�1j�2z�	_��UWM�]^ h0@b�#}:vx�*�z��RڸQ���?;�j��d��[�b1�n*�yL{:�>:mG��S�}s���I���id��Kׯ�� 	`ޫ( ��t$�Vkg�O��SOIy�V�{�*=8��!}$ۘ�g��L�q݊ ��eզ�����ή��ܞ�TJ�-]z�<�� @� ��Y�#[�Cɿ�Ҕ>V%�7���d�{߫�W�j���R���Sߙ��CfYV�Je���ߨ�������YM�aw�Lg�L[o���+V<p��7�H  !t ��x�5����·������~�������\
��������jj�ק��7��>��P�d�#��t�W:I���l!��0�ah��)0q�y���Y�E����ɏ, �:�D�o�g�!���Ֆ�n��X���+����q�2��V]G����(�v�O�ǲ�_ �Ӂ��(��ü�֙��(��i�(���+W^q>�H@[�Z��Z��Ϫ-����7o���
ټ~�t/[�f�}�8�L��@���Q��z�>�����\X����.{���y�������{Z���׭�V  at m#��g-^�Zm��Od�駧���/�(�M�d�?���.m�0Q�Z�˖v�0��TQ���;R.��K����2yJ{]a`��-]z���� I�v?8 t6+���s�tq���.	�S[����{ߓ�NP3?�����kU�w�+K��j�07}J{]};W����o~3/ �@m� ��c����-?����xc�o��g���2���W�˗����L}̡���,���r[�W%aJ{����ͥ7���	 $T[�  ���}�3j���d�=��
�)}<�6}�w��j֟���}}-���w�t�j[#�@3��jqD&Z��{�}���iGI��^71kV�O<I�W  �t mM��>p�)�Y�Pm��v�w���,��7n��SOU���.��:Գ��F�8�۞ڻ ޑ��>��:���=0P;�{���J�8�a���:Γ"p]U8唏�񵯕 ,9�� 0�y�%����~｢GԧJ�������K2�O�De-j����=�2�㨬���HU L;��d��9�،������e�����Oҳf��?��D�d���춝�����[.��w� H8@ǰ]ך��J���P|�7����Аl���Y����\������a�u˲��y��^�(��J !���p��I���?ܵ�אw�g{�;��fϮ�8�u�-i��u;�>���o��S m y�� 0E=�c�,Q��[��qlj�������/H��Wj��N;M�T�������ܹi5oތ�Yg�W��'�,Gccl*�A>��u�q9k�<��堿��Y���_���uW�ƤH⨹V����?���_	 �@Gr<Ϛ��K���j�~4-�]�i��='3��^�}�1�5��Bq�KU�-[֛:�؞��7%��o��Mj�oL'���FFrf�t�ҥ��ҥi�d�Vm����F�͓�_�BTd��I5�B�Q;���/~~ݺ- m"��� 0Mr��֦���/e��G��F�����&���|�>����u�R�,\(�ŋ�L�(᫯J���%��Y�aEQ����,�稣�q�Oz��?�ޠ��S%3��z��Ӳ�f�%uԼn��U?��7�� @!�t<�6}�> =K��Fӫ;vL��-o�R[���z��3B=�$�dD�;N��6���kRٴI��twѢ���]]�a����R�ͩߠ[t�%J�iW��cHҹ��3t�1/��	 � v�.\h-��R5�a��|�ڔ�)SJ��M�h���W�g�����T�:n�"I-^,^�b���-[�S��Fr��={�Ҝ,]�Q}}�{�f�-Ouw[>�鷏b{��}o���:̓r����͝[�,Y.<  �nt ؃�JY3�菤oŊڑl�>;-W��;��S2��sҿr�8�tq��M��k�=����$}���J��z-փ�+��RG��������)բ:���͝��~�������Z��;Y����׬) �! �����{�N8A����6�]�ʏ<�Hm���U����S���������,[&��k|���_���u���,ϳ����%K�j�|7.Sc��Y���fά�Vn��k�0�B�U#���Wq�?# Цt x]K��6�}�	�q��U*��q������2��c���o�z6+�	���]]"˗K��Dv�h�f�n�(A�yF��{zj#�jѢ��Q�G�M]���9�Zx���5kv^z�Lg�-�����S��o�� @#�� ,Ǳ��^�L��g�z�q-���Z�����POuw��j#냃�+�v�,і-���T�x�6�h�8����۲xqV-��̙��I���O��/��C5,Γ�;��l]��ы���� �� IO{_�яJi�f���{�G�t��Qu���}+V�F�ݾ>1Um'�t��f=u��QJB�6I巿���Q�~�牷h�8��y�J�R����0�T�����96�ȵv�ξ��#��z��~v� @ �`����[�W���믫�w�-���i��z�z-ԟxB��K�>Gy�1����vWs�_ݧ�&jxX�8փ�[ŏ/��m8D��I�(_�@��{!����>�\��@X*�����KX.7�s�0�W�Lg��آEc�O?�HٰA �� nb����7��6�u��V�s�S��>+;�wZG�t�N<�|��.\X���;��D܀A�Nz�?���/���##m�.�okG7N�vhKvW����+�q�*���2P��-���ܩ�mzԼQ��n��^�g�.�����ϸ�j�� �:��[��h��7�o��%m&�1����Y�L�<�h�����H���i�����ś=[�N:Iz�;Nlו$�M��Ov{�cr���ھݷ�z�Rݸ1�n��zt�Toomd\_�������愱�ߝ��שX��Wk�`�76�ko�0�JՑO<������#4  !t w�w�����.;v��_�ٱì3ŦI�֌3ΐ�OT�zӷ'���Q3=�~��?�����+�o�Jq��%Itx��g�࠾���*�Td����m���P��ysML$��p��L��C|�,q�G�yoo@(��<L�f�Q����k}��m��� �Ogog����+��ºu� �0:���������K/=���/΍���k���Y����eƙg�����y>�#�z����裏֦���t�d�,I�hZfVe�̜����|y��J)�R	Վ�54T��m�-[�(�'�&��#�ٳŞ1C��3Ŏ�<�㲾�[-��?Ae۶��o�=7���{�0ׂL&�8����v�} �mo����k�}��V�>�~��f
���jxN6k�<�,X��a��ש^~�v�t=���jKu%w%An���o����n|��NP��(�\~;ڷo�:ڷo���q%l@�zzd<�;��!?�ˎ�\��I^r���Y�h�>jq쩧��ysC?W'�����z�_��ڵ7	 t(@S�7^?�#�������L��֑��C��䓕��ڈP���Q��/d�HבGJ�'J��å֨�F��Kǖ9s���E{ZG�����P����h����
v�؈�1��q��Ċ/[_��qGd�Ǜ%�gm��Im���gd��g:Z�uZ�k:·�:�?}����. ��t MG�m�^x��f���g; ҵT.����)�(�z�F���P�/�T�����˥7��3fH;��"�tw��˓��Q�8�=ێ�|>��x���@FG}dD���ؘ�j5�øf{^mD\o�f��j׮ W��{���{d<j��A����?/z}�t��?�暎�g��w�|� �p:������oב>+��L�D��d2����Gf�q���󡇬��lRLL��Cծ�������Ү����pwݔ�i����Y�ʉȍ� ��P�T>X�bǼ��]�s�������J�Ƿ_V:-V6+v�ˉ��8���R�?�#��������@^y�6R^|��R�F�]��g������? �@�::ү��g.���_^�J5d�R�x6}��У�����a�O��՗>�]O}�9�X�:�(��H��F��N�o���A_���q�t �z>~.q�I�Y�J���ڣT*�}W�R�J�W�\�JEſV���M��\W�L�rzzlg`@?��^���{���G[�1�+������G��I�Jg�G�'^x��S�����Z�y�����+�p��`@K]�nݍ��zuiƃ����3����8��U޺Uvơ�#�Q�v�����r:��z��w�KrG!v��$��v���jI����71tTբ>~n����~{����h�CO_:�j��a�k;~�G�k��a�DGZ:]�������q�ڙ���?������G���8����n�5��v]u���}�����_��o~#a�дϭ�\��w2?�����%7�� ���wc ��פ��g>�'�6l�I���+*3w��?�\���^y�Q晆�S��qX����k�u�wsLm���F���y��_���^C�Z_���\ϲ}���4������d�2�;u}���8����7�H��^t F�|ݺ���袳Ԇ�w��tt�}}��R����I��e��':�]ӣ�zzo|��ܒ%ҽtim��+2�$�Ǣ����\_a�����������˅Cg�y��7�p�  � ����Y�ȿ^x�J��c����Ѿ;�$���^+�����#���Xo䨺�G�wO��m�,\X]���Y�0]�ϫz�7n�Vl��4�?T���G�8��?�f�O �O: �\~��/���a���#/��f��F�6���}T[�F�5�����K6���c�+���a�Im}4�bz������Rx�U}fyKv�g�|�
�f��O:��ϭY�  ��@`�������W�����/���B�n{��O���l����L�F���d�'j�]OϞ]����Eb1b�&�GG��T���:̛����0Z���-Y��]��]�M  �@`�_s���^|�?���'�<��?���T��#��&o�G�+[�֮�j��Qu}�/����ǁ���gs�(ׁ�J�~D���v��o�/?����G �A �풟�����gw�~��?�رz���j�ժX���x�3��4'��̂�+�p�d��c���6I)���[oIuǎ�L[�;�OB��jۊ�����N�_�J  �@`��w����?�ڰ�
�Ze����a6u
���n����4}��uo�<��?_��d2�yB� ��А�u��*���b�|���g�)��~�� L
� .���/�ӟ���o�v�Y铡�BO���ꪅ#�z����K_��@I��8�k���T�hoc��?<,�-[���H�A^��\���B������T��h�������|� ��� ��n�ޚ�����<�xN�Gp��4!�k�ϯ������]�-=>=c���̑�5wn�h7��������Q�U��}{-���Vn�?�(g]��+VFW���Ϯ[�1j p�t �r�7��ʚի�o޶�Ł-[x��q'=IF��.z�q�%��]�����*��>n��8sf����@o�7m�w�J��8�+q��_+���`����y�[�-Z~��u; p�t �s�ڵ��aњl��eo����Vi�h�8i�s�HO��]�W^����p��S�࠸z����To�>���,,�����W���^{�Ϥ)���ק���[��X��'~���e� L� �.��ι�3�����z��g:��S��s�`7et��pף��8nK���=�קGߥ�_:���~q����_���E���z3����s��S�'��h�i�}�����
 `Z� ��u���������g}�]�܁O�=�F�3֍�=(��y���}���_q��Tw�8��=����l�vD������Ӽ^��G��|^�BA��һ�����;��_Gժ��z�3u�q�z�U�>��u�� ��!�$��֮}�_��/�O=�̱��u�щ*�u=֣(�g��u�:H�(/�q��X���qqv:��c���_����ka���z���?���>^=j�8ֱ�{��^z���{:�����֣�ah��"\�o��jA��9ߗv��9�䍥ߞ�y�1o�-Z������ ��"�����[�B�]����#{�+�O>���T��G{҃�����Qg�a��ۼy�tZ�X���շ��i 4�����喿��'?y���w�sĪU�n?w�M��`Oʔx��5�f(̜Y=�O^�n� �0:��s�M7=������'���1����;�x��lﵿI[Î�!���,[������]uUQ  E�hK�UW�֧}���������y�c'|��$�{{=҉�ζ�4u������Fç��O�_���� ��t m��o�/k/�t��l8fٲ9م) �Cl�h��B{�3�O��E���˗��%k�<" ��!�����^�1~�w]_߿,ݺ��9'��P���7�J�'#����9�ğ|�G?��<�  ��@�1.Y����r�%��v�=�8f��~o��!�)ܵ����{s��,��3�p���ҥ���7�' �� �t��_wݯ���]]7����u�)��8�E�k�|]=������o�
�=���F͟|R  �C��H����O��E�0p�}?;v��Y�E���6r0Q�������~�d{����#:������˖�Ǩ9 ��@б._���a�����^��k��;��r]J�CL6N�����Ow�����������6F�NG�W���;�8O�~Z  f �t�o���5���?�x����>��YFӱ{�/!�D��qĶ��G����_��  �B�@��|��a�.�ે���Y|���TO�m����+����JΪ@����:{w !�@� ��sʨ��TTF8#;�g�IUu'3�m�򠻪9�9Td�ħ��qDf�����:.@P���;�T�[�փʖ�Iߪ��ι�ޯ�!��!!�|_}������<�v[  =�1.\�������Æ:*�{���(d��P�V�������>�`�+�y��[ �� �e�W���5מwމ|�Y�d�ܙ�.ҁ�������g��n�r  y�	�s�շ�i�U����E����>���:f��@򆺺F}�����O}jY��7 �A�<�w�[�7k/����6|����_;��uv:���i�j��7�8�ug{���t��a����]w��6�v�-K������;Ϋ��$�����G���E�\|� MI�솳?��{�t�u�{��/}��#=�G!ҁ��86��~�s�;��k�) ��:�8��k�1N�?z�2�k_���gwM;�@��3�<pp��ǿ��O|��� @�� ���7��8}���O��E��_���?�c���:��Ξ=���n8�3�9?l�4;@+� �u��[��}ߵ��~��o[p�1�Y��:0a�b�o>���{�ao?�� h9`�d}}�8�=�z�;������3:��)��B�c;f��|�1_�w��o;K��4�0��C��u��v�}w����ccg.��nzl��#�ڂ@�KN_�~,N�X{�K����?�(�S�:�T�ۯ�(�M;,8s��G ڄ@�������ƣ����+�rgt��:f����m�3gx�s�s���g	s��$����G�/h��N;��j����wN?�� ���c��G��N����' hS`��~�����'��÷/�ַ����:�,��:��Z>=��?���}��m�v֧> ho`Λ~�϶o�#����
Y�ߞ��L�V{�#~6�x�;ξ�����n �+����Y���O8!�7:���'���p�a��|�:��g��r��_�-��3���  �C�$���~y���q=����4>gN��hQ �K-��.ܼ�#n<���.��r ��@H����Gq�d��p�~s�,	�3������MK��9|�A�������O~2 �S� �k<����c��Z-�w�]a�#���1ܳ\. i��_�[-ڴ��C?6#�_~���c v�@h1 6qĮ�;¼��$�j<��iS &��Y�F7/Y�!�x�Eo���[÷� `O	t�&4<sf��B�c�}������0��?��� �]cS�ֶz�C�]s�1���ϖ0Q:@��~����'���+������4dc����2�˅mlٹx��p���~�54�~N ��#�ZD-���,�5��?�a�ڰ!�ݸ1�C7�`�eY�6o���!�|;7oޟ���>���� �[:@�:5<z�	��/�l	]w��k�/~B��'�|�ܹC�/�04g��w�[��!���}A����ٳ��/}�1}ǎ0#�z�����C��:�z#���ܱp������Y7�pS�� �k��͜�����)�_�X�2�G?
��󐍎h������ڲ㠃���?�笫��ݝr &�@hS�7�?��1�g����������)��Zͮ��|�#;.�%?wn錫��/ @B: a��#l>�]��Z-t>�@��яBW��·
u��ӄ�]ڱ`�O�x����˧�;�7�  E�ߐ�r�>���zU�24�6n3~��0;�ԭ[�jdƌ��<�}��[k�g���7�{t�&!�xR#ӧ�G�����y����C���u�ݡ��?��;L��ԩ����oZ��?��s?p�7��� �	t v��y��C/yɮG�gn��� ���8�}~��h�ap���}��)S�\��ғ/��t ���k<?x��F����`����a�ƍaz���fl���^gdY��?l[�0�8䐰c��3^���X,�/ @� L�F��?�/x���Mٱ#L���03�Y7��|�|~t4�[ƦO�<0�xֳ�ТE��|l֬  �B��W�̜F�:*l��^�_V*����s�9)�u���M�^<�G���ó:��E{������A�zd}(�;��i�6 Ю: ���^��8}�W�ߺ��)�o�|f��Л:6o>nʣ�.���3����<��OUuu���s�Ё�
�F�Ϟ ��$��t/��ʑ8]=>~�K�.|xӦ�;�m{Un˖%Ӷn�;m˖S�o�Ȅ{Z��0��~���cx��0�x���9�>eJ  ��@ YoZ��q��ߌ�_�詧��������m�߱�)[�ԱeKW�iS��}�wt����a��ٻ���!�3��P��F� {N��tο�G�t���7�u֬Cxmmh����O�28�8F��8��ǀ�>4��FF|��q4�t͚����{��q�Zϙ��3���G��RN��Ƕ����������ux���Ν/��G憆���?�s笸��1<<5?4�1m��\nt4׬��5�)�M��bX�Μ�k�� ���a4εF�7��Qt �T���k��+N�q�S��[O;m�]�����gg��!c�Ë���룣󲑑��cc����N���2�)cc����)Sj�ldl�#�=S��~}�9��ƗBG�Z-�?��,�5�6����\-�kYVi\g�X.���8������)�cC��S����cӦ�<�SkӦ����?���xI �: <�ׯ�ӆ�U�VT��N��{ ��@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@ �N�^� ��t ��dY6�\.�*�J� �� 4�\.w\�� �Et �)�j�7�@� @Sʲ��8�? @�� @�z^�Ryy�X�j � ���U��q� �� 4�,����������� hr ����h=�˅6����z�����  ML�@���>2u��Юb���Z���� hb ���ٳw�vV�ׯX�j��/_~ �&%���=���C����,
m*~�����>C��u�Y	t hr}}}��J�Ѹ��X�7�}�(.� hB Z@�^0j[��U1ҿ�lt ��@����8�\܇)�z��+����y�{~ ��t hw��@#����~����5}}}; 4	� - F���w�=�˺����H���g� 4� - ����o;%F�Uqo��fw ��@�022�aʔ)��qv�R�+�� �8� -`�ʕ�����,�~Cܓ���~�X��  	� �:�%����^��Z�>T(� H�@��e��@\qo�Z��Jej�X�> @�: ��[�ő��F����k��r�T*]  1 ZD�X|�R��G\�0��#���j5+
� H�@����1B������A��� ��8�"�~u'�\.�K��G $@�@��yG���b��4�T���H�R9�X,V L2� -�^�_%П��OY��1��
��� `�t h13g������������Z�.�����o4 �$� �b.���m�r������ܮh���g,[�lg �}L�@���Z�vNp&��z�����c��#}K �}H�@Z�|��J��ٸ<5��^5<<�����7���� `� Т����*�˽y�Eh솸e�����8����� �� -����;�r��|]`O���\�TN+�7 ��: ��,��:�g�+���HG��� �E ZX��[c\~:.��SS���u�r�٥R�� �� -ntt�='�����o�R9���ki4 `�	t hq+V��'�e%.�x��߲eˢիW��c� �h �@�e�5�E��a�g$��kGFF�r�e���bŊ{ L� m�P(���R\�L��vtt|5��J�� &�@�6C�J�Sq���D84˲��=}s�X�j �gH�@{YZ��/��aN��.��g5�$ �3 ����Ň*�ʅqyS`BdY6-F���j��B��6 �� �fb�&F�uqyv`B�H��H�������] `t hC�|��ccc���&RO�\�ܶmۻ���j v�@�6t�%�<Z�VO��j_n<��0q?/���:������ �&� m�P(|�\.������1�s1��� <] �X�TZS�T^|}o8��k׮=c�ҥ# ��@�6W���4˲�屁��G[�n��z��-[�lg �'!��͕J��J�m1ԿC}��D;eddd}���D: OF� ���~P.���7�150��4<<�����m>��� �.�R�K1��,˲&\��7wvv^#�G��x: �k1�?#����.��]]]��z��q] � �۶m+ň\��������8_ �1: ��_���3�,�%^�,�7��R�<X,�w �q ��7�W��7���������-�ˏĽ��  A� O�P(<���r>��j�<<�7������� @�� ����/�ks�\#�&T�e�8n(�˯.�J� hk xR���?�T*o���_�1�`�͌���_~��.�䒻 mK� O�X,�G������/�&ڂ����]z饿�r��M��$�������;��r���eW`BeYv̔)S�a���'-[�lg ��t �i����z�Ry]\~>�������W��� @�� �n)���>˲����PqO�)���^*�> h+ �m���_���z��Y��W\���{OO�W mC� {�T*}�q<X��Ɲ���	�sJ.�[_�T^\,7 ڂ@ �X��oƈ|M��/Ĩ��0q?������ޗ���� �<� <#�#ت��k��-��L�������j|�� @�� �3V(n������s�&ҹ�r�+�R�#��&��	������/ϲ�qN�с	�t����7����3 в: 0aJ����j��Z��x�����2=�����/�yt��%��	U()��'���8^�1Џ���"./ �$� L�R������;;;��a���D��J��o�b�� @�� �^���7#��鿌��,0!���n����I ��t `���^��{*���bX^C=<#qg�qݺu�^q�駏 Z�@ ��b���Z�n���8*̟?����}���s5 �2� �'
�µ�ryS\~"˲�g�oW�Z���˗o �� �3�R��j���z����{,˲i�Z�ڵk׾t�ҥ#��'��}�P(ܶjժߏq������3�[����� MO� �\�������|#ҟ�c�z�}�j���B�� @S� �����o͚5��1^��#�G�/����}��[�hR �4_|�u�֝z�=�����
�Ϛ5�q�P �i	t `R������J��J�sq�.+��7�J�_ ��@ ���w��vK��q����� @S� @2��J�7.�o�����j�zm�� 4� $�T*}qժU/��j�������������k�>��� �G� �i�V�VOl����vǱ�7o�(�W ��@ �T(~�z��W������'��\.���/���K.��� @�� @��-[���������5Y�-<]�����sO �it  i}}}�qzW�\�Y�/u�����q�>X*�� 4� 4���18h��sJ�L��o�8; �: �4b�_300p�O�ˮ����tF��===�	 $O� M�����j�5�z�q��'������� @�: �t
��7.���W���ޒe����9�R��X,o $M� M�K.�3F���#������7��) �4� 4��w�"������獕J��b���d	t ��uww?p饗�����s1D_x\�w��( �,� 4��+Wn���?)��5"�����-�V�:n��� I� @K����#�1�?c���oˍ���E�� $I� -��W�~�����w�]qON��˺W�Xqo  9 h)˖-�#�u�����cu������ @r: �rV�X�9F��1F��e�K���իW��e�v �"���4�'utt�/_�%˲�###���_ H�@ ZV#ҫ����������~� ��#���V(Y�z�I���_Ͳ�@��V�Z���˗+ �� ��e˖=X�VO���_������q� 	� @[(
?xm.��r��/��,�N���}w__�p  	 h����Y�V�R���)����tvv��� � ���R(��\.���%i����  h;�R���s�,�?�������.�l���� �N� m)F�+��qY�kz>���8_ �t h[[�n����zN\���ۃ@H�@ �V___������|��xy|hCY����5k:/���m�I%�����ӳ�\.�9.�cu^h?S� xY��� @�+�J?�T*g���B{����A�L:� �ś���_gY��L��_ �t `ܶm������1XO�������{zz~ �4 `\�q�W�>{dd�����F�,k<�.�&�@ x�e˖=X�TΫ��7�h�B���r����I#� ~K�X��\.0./
m�^��$ 0�: ��ضm[wWW�k�����,;��.[�bŊ{ �B� <��������vy�=�˽8N`�t �'�����J�rU\�3���@�t `Rt �'�eYw�V{s���s� �K� <�B��H�R���PhqY��  0i: �S8�C>z��w/�{Lhms�����_J �9� �N?���r�����Dhq�z��8	t�I � ��b���Z������e�q�v `��  OC�z�\^�kC���$�  O�ԩS�W[���`�t ��iٲe;���5qY-�t��#� vC�e7����� L
� �
��w���q� ��Y�I!� vC�eq�J�qyFhM`�t ��T���=�zKz�޺ �B�L�����-��'����5�Z�;� �D�L�+Vl����t�,k�@��۴�k�NY�t�H `��  ��X,��l_��k֬�ܺu딽��\xᅣ1� ��@ h_|�}��\�2 ��	t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H��@\��@PD    IEND�B`�PK
     `_[�kZ��  �  /   images/6608fa58-7afa-4488-b64c-2b761d69d6bd.png�PNG

   IHDR   d   }   T;�   	pHYs     ��  �IDATx��	�U�ǿ��ʪ>�/�FA��V�i<vD@YqWCא��Y�q�Й1�u��	cw5vv����@Ggt=wW�G%D9�� ���>��:�z�}�UM�4ts��������ʪ�z����/*%��@$S�d*�LE ��D2�H�"�T"��@$S�d*�LE ��D2�H�"�T"��@$S�d@v,X ������u�a�y�3!��sp����C�\��0�$-�P�������	���ǡ��2�YV0V�JqS�-��;]���jl���i��l:�L���*8g�z�����A8�pǁj�PUu��
���bg��Q���ld&.6S8NW˅~�p>ö��5�̄L��i�S^6n�%���f��ɓ!���0����_�����\|���wr����(AQT>��G���H"���5l/ۺޮ �C]�ee0���@FI��W_�h	.��:aiZ=��?������'�
��+�m(�(
�;�<�V��<��7��{��&���`綾��@6Ȏy󠼵���cS}���m߇o�`�b���Ex�+'��)��{��8�@:m��Zfs�����5�~����?{6�ߴ	dRA��x�����t�������=-ŷ2^C��\&5�lV���!jn{�koݚ�7o6E"a���h-W���OWQ~�ZW�~g]|��;["(�u�"(9xЃa�j9�U�a�R�x�C(�Q!	�!8����J�WTp��!��Յ̵k���m�/�4Y���b��?�ٽ�Ν%��
���҆*��Yy�ʤI�~商��Y��O�L�Nl*dI�	�G��ٳ�|�X�
�����Q>n\�\��a�D0%��>�Pno>��MQ��_uL��(�
����]���R۟#�� ö�6kVH�??���,W܎��� �A!k۾ݴw�/Եy�f��M��0/)�w�I"p��2���Sn��`�2(p ��.�ҝ;�MA��d��� �A�K/#Ë�7B���̫�&�x�����;PUF�%�rZZ��u�EYY��R�?_�%堘Hw"Ɣ�Fm���0��ud̡C��؀���џB��@7�Μ�!�L��n�P%�dI4��	�J�A=��к������o'�˖���C����Q\��%�ֹ������l�5�NC�8�/�L��E��{�3&�*�t>f��/X`x�a�u2��L��f^��&'���	�k1��LF���ffv?ʆ����v���.�Ik�B�(���c�u���Ơ���:���+�x����qج?�)c�Y�F+�=)aǻ�9���yO�)�i.C0/�`^H
����\�Xk`'���ۧMө�;
����}Xy�4���;����4~�����(���D��;�d�=��"�Ǥ�!*�����k������I�� ��c�?����5k�
Ⱥ%K@mj�[�yf���)v��(��*��h	��ۡ�"ﶾeѾ#h%�s��|4&�R`@�����t�������UaFt����[��.�A�3'O����WWC��DY�w�I06��r��=��+��lֵw�0���\�9�55L8RP $��*Z���x A�-}����wWT�S;� ~jr�B*�6�����  ���6fL%�7�#*Ԏ�����r�P����D�ߝ�)0 X	��f�4�[���A�+��m������:P����)/�*|�^�	�c��}�uM�چAz*�T�K�A��)<E>ӓLR����~&�+��<�:�qL�87��E�!�uZ��X�ǣ���\���7�.K���0�
<S�Ϥ��1�pg:j����)���jBUU��� �Ud	���*'9�0����T6q8W���)�ӾaT�z���t)Ĳ��Bb �� B�����8
���4�,��n*U�F�㔠�U��%�� ҫ�Lw	��ya�Q��oK8N$n�U0L$����1
ap�:=$1^��f�;�*�$�
���鵴ㄆ҈ p��Lg2�S.˹w�k���4�`���������EuSҊR���p�A�@Y�"�EnK0�3��i8a��R�0�𣆖C��o��9���B���s\�H�=���}-�K"���	��ؐ.��{c�LF-	�L�/�k�bY��1e
���W�
<ǎT�BP�T�u�s]��{���ڜ�����k�
2�Rð�
����o��f궽�v�xv�,�~c#���33m���,�5�4���I�	&9�>�Љoy�FxӜ�;�G���w2t�RzY$b�"z����0�����[*��U �CI��J�ٱ���;u2�y(����e"��
�m�뎋:�ӟ�xc�w��G���3a��_BP
���?�MP'��Y�����1�h)d�]�۵L�u�]����y����x�3w{�x�Π3n�ݧR��a�Ŷ��]W���{�Z��ر
�#�sf���ꄂNj�/ʼ���=G0�̜�c�\�k�}�l�+�CB�J=�N*9�rA^��]�q�R-k͝㮀�#0 6����g6P(2�H���3M	�cfc�uu [�@
q��(�e^ַ�A�{'���Ye�f.�H�������E�t�.��P8'_f3E���!N����I,ӹ�W�q��w]�9�Ht�tP
H<��V� �g�:�Y�ug�;�[�D����"�p}�����bY4�A)0 =�ࡇ ��Sj)�u��x/ZB��P(��#���}��Gi�;�%�δe�Wsy~�>�U�io�]w�h-kۚ�(4(rUx��{:�sΦ��� �S	�6Z�)e��l4l=��@K�٬�����^J�!Ť5�����@�(�y�)ӄ]���Bt<��(�����h~��ؾ��2�KK;��IOԆ�R�L�̿�� ƒ[����R�4I/;
��*��H� �	��Exh,-��3��r[�2:�pVd4#�aP0��h�0�fiG��w�~J��cG �UU��^S^���,����%m���i��Y�Q[�ɲ�mCɥ�?�7�o�W�\ ����uYc�Q�����}�Z�::��E�X*Y�2�P�T��"pr��'�Ώ�>G7DIE�#�.�j�ca�u�h��][Z*�r��BD}�:u��ܷ��Z%F-\�J�;O�3%����_�����������pnG��ŪT��ٶC+	��h�e��H��)T�7f�>��P�'������K��w킠�T=���a�;[��bU@ۚ5��[o	�t��3Q[��	J�%K"��_���2��Np����c-�!�*�����KU�����	a>u�a�b���{�ݸQh�*%��?JWQ6���>d��C)���<�$��w���������D��d�5�l���]+�^~��&b�fqc�d�>ܞ--%X�"�EO-�*h)A�q�������%:���~��jZG�)��1�`��A����=��E��
 W��WV4zS��9M��<k�HB�E�0�:w���TV�H���p7�%���.]��x:6n���^;42iD�9Bc�j�	u"so�9ArmD�4N+C@n���Hߗ��K��%2MM��k
&�v̀Ch[�R5�ٯ�&��+�@�
H�5�@����)S��k��Ic{�l����ara�1��3��7���م�;T�D��g��3��L--e
Z�7I�������$�]]`b݀	8�8/��m�p��a�7������;�D"N0�'O��?�
���,�Yx�?��իa�����{�Y���7E�����\/&�AA�
>��9�N��--`�Ҳ�U�c}��Wn�k*��c!x�y�a<:������:Yta,��.�h�u�ʕ��'w��y�>��g/��g�����w��c��s<���{��π|X���z�6�_�=={>�:�2��n���*�Ĩy�����	gc�Xtｎ�l߾���ӧ�_0�V���)�ӹ�з�#S�9?��'Zi��[)�-A��5
��J|�^(�
6S�W_�?���5����:5qH�ZU�#�[o���;�t�c,�9�޲~��{�:4�E�E�ob�~/��҆n
Z������믇�o����S�\�
�x�	hŴX�ʙ�#y�Y�8�l��tҕ_|���u�c�!�����She!�|���Ucq���b6�����A�׎jl��"T1M���`�����u�OkS��$
���,��ĈŋW����aG.�L�/�8����$������[�lT�����̯�us�Y���zOj�88��� ��W<����m�@FI	�W9�%�����8x�F zg'�,B��CsC���"13'%��䢮�Ј��Hn �t㧟����G�+d�&|�V@�?�D2�t �ʼO��< �k� 0��!l�`�9�1�� ��Z��$���(��*Q١{ 4����Z����lB.�E��g�����a����l�@�U�
���j،~�o����O�7FB{ ބ6�������6r�?�?���!���@V�X�ulN�`�۪|��Ѥ�_H٠{ $��>P��?-&(��}��m3ZWa/~������/�o��؜���fc��JFR?(侮��_��`s�ӀҬ_0��VQ@H���F~�����b{�?������B�5‐�A�3����!�(E^��%Y�D6 �F?���|���=7��dA/�$�ݦD�D��k4���K�����
�ŧc3��Uh�kH$)��0=�;����@���ө~w
󗏽[i��� �]\}%�>����C�&�� �m� < ��ȉ$����D2�H�"�T"��@$S�d*�LE ��D2�H�"�T"��@$S�d*�L�I�����\�    IEND�B`�PK 
     `_[�X�,�  ,�                   cirkitFile.jsonPK 
     `_[                        Y�  jsons/PK 
     `_[1G��  �               }�  jsons/user_defined.jsonPK 
     `_[                        ��  images/PK 
     `_[�R�W�  W�  /             ї  images/e30496d1-6e1c-40fa-a66f-2add70ecdc94.pngPK 
     `_[$7h�!  �!  /             uB images/a7fde0f7-2836-4f0c-aad0-66dcccec46ff.pngPK 
     `_[wJ���  ��  /             �d images/f9728bc6-2422-4ead-9082-90351081a874.pngPK 
     `_[	^�G�  �  /             � images/9ba3df0f-d630-43f7-8169-617793654d93.pngPK 
     `_[�e�e�  �  /             � images/3d0a314b-f708-4b2c-819f-35c414b123ec.pngPK 
     `_[�kZ��  �  /             �� images/6608fa58-7afa-4488-b64c-2b761d69d6bd.pngPK    
 
   >�   